/*
Copyright (c) 2019 Alibaba Group Holding Limited

Permission is hereby granted, free of charge, to any person obtaining a copy of this software and associated documentation files (the "Software"), to deal in the Software without restriction, including without limitation the rights to use, copy, modify, merge, publish, distribute, sublicense, and/or sell copies of the Software, and to permit persons to whom the Software is furnished to do so, subject to the following conditions:

The above copyright notice and this permission notice shall be included in all copies or substantial portions of the Software.

THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE SOFTWARE.

*/
module afifo_35x2 (wr_clk,
                   wr_reset_n,
                   wr_en,
                   wr_data,
                   wr_full,                 
                   wr_afull,                
                   rd_clk,
                   rd_reset_n,
                   rd_en,
                   rd_empty,                
                   rd_aempty,               
                   rd_data);
   parameter W = 35;
   parameter DP = 2;
   parameter WR_FAST = 1'b0;
   parameter RD_FAST = 1'b1;
   parameter AW = (DP == 2)   ? 1 : 
				  (DP == 4)   ? 2 :
                  (DP == 8)   ? 3 :
                  (DP == 16)  ? 4 :
                  (DP == 32)  ? 5 :
                  (DP == 64)  ? 6 :
                  (DP == 128) ? 7 :
                  (DP == 256) ? 8 : 0;
   output [W-1 : 0]  rd_data;
   input [W-1 : 0]   wr_data;
   input             wr_clk, wr_reset_n, wr_en, rd_clk, rd_reset_n,
                     rd_en;
   output            wr_full, rd_empty;
   output            wr_afull, rd_aempty;       
   reg [W-1 : 0]    mem[DP-1 : 0];
   /*********************** write side ************************/
   reg [AW:0] sync_rd_ptr_0, sync_rd_ptr_1; 
   wire [AW:0] sync_rd_ptr;
   reg [AW:0] wr_ptr, grey_wr_ptr;
   reg [AW:0] grey_rd_ptr;
   reg full_q;
   wire full_c;
   wire afull_c;
   wire [AW:0] wr_ptr_inc = wr_ptr + 1'b1;
   wire [AW:0] wr_cnt = get_cnt(wr_ptr, sync_rd_ptr);
   assign full_c  = (wr_cnt == DP) ? 1'b1 : 1'b0;
   assign afull_c = (wr_cnt == DP-1) ? 1'b1 : 1'b0;
   always @(posedge wr_clk or negedge wr_reset_n) begin
	if (!wr_reset_n) begin
		wr_ptr <= 0;
		grey_wr_ptr <= 0;
		full_q <= 0;	
	end
	else if (wr_en) begin
		wr_ptr <= wr_ptr_inc;
		grey_wr_ptr <= bin2grey(wr_ptr_inc);
		if (wr_cnt == (DP-1)) begin
			full_q <= 1'b1;
		end
	end
	else begin
	    	if (full_q && (wr_cnt<DP)) begin
			full_q <= 1'b0;
	     	end
	end
    end
    assign wr_full  = (WR_FAST == 1) ? full_c : full_q;
    assign wr_afull = afull_c;
    always @(posedge wr_clk) begin
	if (wr_en) begin
		mem[wr_ptr[AW-1:0]] <= wr_data;
	end
    end
    always @(posedge wr_clk or negedge wr_reset_n) begin
	if (!wr_reset_n) begin
		sync_rd_ptr_0 <= 0;
		sync_rd_ptr_1 <= 0;
	end
	else begin
		sync_rd_ptr_0 <= grey_rd_ptr;		
		sync_rd_ptr_1 <= sync_rd_ptr_0;
	end
    end
    assign sync_rd_ptr = grey2bin(sync_rd_ptr_1);
   /************************ read side *****************************/
   reg [AW:0] sync_wr_ptr_0, sync_wr_ptr_1; 
   wire [AW:0] sync_wr_ptr;
   reg [AW:0] rd_ptr;
   reg empty_q;
   wire empty_c;
   wire aempty_c;
   wire [AW:0] rd_ptr_inc = rd_ptr + 1'b1;
   wire [AW:0] rd_cnt = get_cnt(sync_wr_ptr, rd_ptr);
   assign empty_c  = (rd_cnt == 0) ? 1'b1 : 1'b0;
   assign aempty_c = (rd_cnt == 1) ? 1'b1 : 1'b0;
   always @(posedge rd_clk or negedge rd_reset_n) begin
      if (!rd_reset_n) begin
         rd_ptr <= 0;
		 grey_rd_ptr <= 0;
		 empty_q <= 1'b1;
      end
      else begin
         if (rd_en) begin
            rd_ptr <= rd_ptr_inc;
            grey_rd_ptr <= bin2grey(rd_ptr_inc);
            if (rd_cnt==1) begin
               empty_q <= 1'b1;
            end
         end
         else begin
            if (empty_q && (rd_cnt!=0)) begin
				empty_q <= 1'b0;
			end
         end
       end
    end
    assign rd_empty  = (RD_FAST == 1) ? empty_c : empty_q;
    assign rd_aempty = aempty_c;
    reg [W-1 : 0]  rd_data_q;
   wire [W-1 : 0] rd_data_c = mem[rd_ptr[AW-1:0]];
   always @(posedge rd_clk) begin
	rd_data_q <= rd_data_c;
   end
   assign rd_data  = (RD_FAST == 1) ? rd_data_c : rd_data_q;
    always @(posedge rd_clk or negedge rd_reset_n) begin
	if (!rd_reset_n) begin
	   sync_wr_ptr_0 <= 0;
	   sync_wr_ptr_1 <= 0;
	end
	else begin
	   sync_wr_ptr_0 <= grey_wr_ptr;		
	   sync_wr_ptr_1 <= sync_wr_ptr_0;
	end
    end
    assign sync_wr_ptr = grey2bin(sync_wr_ptr_1);
/************************ functions ******************************/
function [AW:0] bin2grey;
input [AW:0] bin;
reg [8:0] bin_8;
reg [8:0] grey_8;
begin
	bin_8 = bin;
	grey_8[1:0] = do_grey(bin_8[2:0]);
	grey_8[3:2] = do_grey(bin_8[4:2]);
	grey_8[5:4] = do_grey(bin_8[6:4]);
	grey_8[7:6] = do_grey(bin_8[8:6]);
	grey_8[8] = bin_8[8];
	bin2grey = grey_8;
end
endfunction
function [AW:0] grey2bin;
input [AW:0] grey;
reg [8:0] grey_8;
reg [8:0] bin_8;
begin
	grey_8 = grey;
	bin_8[8] = grey_8[8];
	bin_8[7:6] = do_bin({bin_8[8], grey_8[7:6]});
	bin_8[5:4] = do_bin({bin_8[6], grey_8[5:4]});
	bin_8[3:2] = do_bin({bin_8[4], grey_8[3:2]});
	bin_8[1:0] = do_bin({bin_8[2], grey_8[1:0]});
	grey2bin = bin_8;
end
endfunction
function [1:0] do_grey;
input [2:0] bin;
begin
	if (bin[2]) begin  
		case (bin[1:0]) 
			2'b00: do_grey = 2'b10;
			2'b01: do_grey = 2'b11;
			2'b10: do_grey = 2'b01;
			2'b11: do_grey = 2'b00;
		endcase
	end
	else begin
		case (bin[1:0]) 
			2'b00: do_grey = 2'b00;
			2'b01: do_grey = 2'b01;
			2'b10: do_grey = 2'b11;
			2'b11: do_grey = 2'b10;
		endcase
	end
end
endfunction
function [1:0] do_bin;
input [2:0] grey;
begin
	if (grey[2]) begin	
		case (grey[1:0])
			2'b10: do_bin = 2'b00;
			2'b11: do_bin = 2'b01;
			2'b01: do_bin = 2'b10;
			2'b00: do_bin = 2'b11;
		endcase
	end
	else begin
		case (grey[1:0])
			2'b00: do_bin = 2'b00;
			2'b01: do_bin = 2'b01;
			2'b11: do_bin = 2'b10;
			2'b10: do_bin = 2'b11;
		endcase
	end
end
endfunction
function [AW:0] get_cnt;
input [AW:0] wr_ptr, rd_ptr;
begin
	if (wr_ptr >= rd_ptr) begin
		get_cnt = (wr_ptr - rd_ptr);	
	end
	else begin
		get_cnt = DP*2 - (rd_ptr - wr_ptr);
	end
end
endfunction
// synopsys translate_off
always @(posedge wr_clk) begin
   if (wr_en && wr_full) begin
      $display($time, "%m Error! afifo overflow!");
      $stop;
   end
end
always @(posedge rd_clk) begin
   if (rd_en && rd_empty) begin
      $display($time, "%m error! afifo underflow!");
      $stop;
   end
end
// synopsys translate_on
endmodule
module afifo_77x2 (wr_clk,
                   wr_reset_n,
                   wr_en,
                   wr_data,
                   wr_full,                 
                   wr_afull,                
                   rd_clk,
                   rd_reset_n,
                   rd_en,
                   rd_empty,                
                   rd_aempty,               
                   rd_data);
   parameter W = 77;
   parameter DP = 2;
   parameter WR_FAST = 1'b0;
   parameter RD_FAST = 1'b1;
   parameter AW = (DP == 2)   ? 1 : 
	          (DP == 4)   ? 2 :
                  (DP == 8)   ? 3 :
                  (DP == 16)  ? 4 :
                  (DP == 32)  ? 5 :
                  (DP == 64)  ? 6 :
                  (DP == 128) ? 7 :
                  (DP == 256) ? 8 : 0;
   output [W-1 : 0]  rd_data;
   input [W-1 : 0]   wr_data;
   input             wr_clk, wr_reset_n, wr_en, rd_clk, rd_reset_n,
                     rd_en;
   output            wr_full, rd_empty;
   output            wr_afull, rd_aempty;       
   reg [W-1 : 0]    mem[DP-1 : 0];
   /*********************** write side ************************/
   reg [AW:0] sync_rd_ptr_0, sync_rd_ptr_1; 
   wire [AW:0] sync_rd_ptr;
   reg [AW:0] wr_ptr, grey_wr_ptr;
   reg [AW:0] grey_rd_ptr;
   reg full_q;
   wire full_c;
   wire afull_c;
   wire [AW:0] wr_ptr_inc = wr_ptr + 1'b1;
   wire [AW:0] wr_cnt = get_cnt(wr_ptr, sync_rd_ptr);
   assign full_c  = (wr_cnt == DP) ? 1'b1 : 1'b0;
   assign afull_c = (wr_cnt == DP-1) ? 1'b1 : 1'b0;
   always @(posedge wr_clk or negedge wr_reset_n) begin
	if (!wr_reset_n) begin
		wr_ptr <= 0;
		grey_wr_ptr <= 0;
		full_q <= 0;	
	end
	else if (wr_en) begin
		wr_ptr <= wr_ptr_inc;
		grey_wr_ptr <= bin2grey(wr_ptr_inc);
		if (wr_cnt == (DP-1)) begin
			full_q <= 1'b1;
		end
	end
	else begin
	    	if (full_q && (wr_cnt<DP)) begin
			full_q <= 1'b0;
	     	end
	end
    end
    assign wr_full  = (WR_FAST == 1) ? full_c : full_q;
    assign wr_afull = afull_c;
    always @(posedge wr_clk) begin
	if (wr_en) begin
		mem[wr_ptr[AW-1:0]] <= wr_data;
	end
    end
    always @(posedge wr_clk or negedge wr_reset_n) begin
	if (!wr_reset_n) begin
		sync_rd_ptr_0 <= 0;
		sync_rd_ptr_1 <= 0;
	end
	else begin
		sync_rd_ptr_0 <= grey_rd_ptr;		
		sync_rd_ptr_1 <= sync_rd_ptr_0;
	end
    end
    assign sync_rd_ptr = grey2bin(sync_rd_ptr_1);
   /************************ read side *****************************/
   reg [AW:0] sync_wr_ptr_0, sync_wr_ptr_1; 
   wire [AW:0] sync_wr_ptr;
   reg [AW:0] rd_ptr;
   reg empty_q;
   wire empty_c;
   wire aempty_c;
   wire [AW:0] rd_ptr_inc = rd_ptr + 1'b1;
   wire [AW:0] rd_cnt = get_cnt(sync_wr_ptr, rd_ptr);
   assign empty_c  = (rd_cnt == 0) ? 1'b1 : 1'b0;
   assign aempty_c = (rd_cnt == 1) ? 1'b1 : 1'b0;
   always @(posedge rd_clk or negedge rd_reset_n) begin
      if (!rd_reset_n) begin
         rd_ptr <= 0;
		 grey_rd_ptr <= 0;
		 empty_q <= 1'b1;
      end
      else begin
         if (rd_en) begin
            rd_ptr <= rd_ptr_inc;
            grey_rd_ptr <= bin2grey(rd_ptr_inc);
            if (rd_cnt==1) begin
               empty_q <= 1'b1;
            end
         end
         else begin
            if (empty_q && (rd_cnt!=0)) begin
				empty_q <= 1'b0;
			end
         end
       end
    end
    assign rd_empty  = (RD_FAST == 1) ? empty_c : empty_q;
    assign rd_aempty = aempty_c;
    reg [W-1 : 0]  rd_data_q;
   wire [W-1 : 0] rd_data_c = mem[rd_ptr[AW-1:0]];
   always @(posedge rd_clk) begin
	rd_data_q <= rd_data_c;
   end
   assign rd_data  = (RD_FAST == 1) ? rd_data_c : rd_data_q;
    always @(posedge rd_clk or negedge rd_reset_n) begin
	if (!rd_reset_n) begin
	   sync_wr_ptr_0 <= 0;
	   sync_wr_ptr_1 <= 0;
	end
	else begin
	   sync_wr_ptr_0 <= grey_wr_ptr;		
	   sync_wr_ptr_1 <= sync_wr_ptr_0;
	end
    end
    assign sync_wr_ptr = grey2bin(sync_wr_ptr_1);
/************************ functions ******************************/
function [AW:0] bin2grey;
input [AW:0] bin;
reg [8:0] bin_8;
reg [8:0] grey_8;
begin
	bin_8 = bin;
	grey_8[1:0] = do_grey(bin_8[2:0]);
	grey_8[3:2] = do_grey(bin_8[4:2]);
	grey_8[5:4] = do_grey(bin_8[6:4]);
	grey_8[7:6] = do_grey(bin_8[8:6]);
	grey_8[8] = bin_8[8];
	bin2grey = grey_8;
end
endfunction
function [AW:0] grey2bin;
input [AW:0] grey;
reg [8:0] grey_8;
reg [8:0] bin_8;
begin
	grey_8 = grey;
	bin_8[8] = grey_8[8];
	bin_8[7:6] = do_bin({bin_8[8], grey_8[7:6]});
	bin_8[5:4] = do_bin({bin_8[6], grey_8[5:4]});
	bin_8[3:2] = do_bin({bin_8[4], grey_8[3:2]});
	bin_8[1:0] = do_bin({bin_8[2], grey_8[1:0]});
	grey2bin = bin_8;
end
endfunction
function [1:0] do_grey;
input [2:0] bin;
begin
	if (bin[2]) begin  
		case (bin[1:0]) 
			2'b00: do_grey = 2'b10;
			2'b01: do_grey = 2'b11;
			2'b10: do_grey = 2'b01;
			2'b11: do_grey = 2'b00;
		endcase
	end
	else begin
		case (bin[1:0]) 
			2'b00: do_grey = 2'b00;
			2'b01: do_grey = 2'b01;
			2'b10: do_grey = 2'b11;
			2'b11: do_grey = 2'b10;
		endcase
	end
end
endfunction
function [1:0] do_bin;
input [2:0] grey;
begin
	if (grey[2]) begin	
		case (grey[1:0])
			2'b10: do_bin = 2'b00;
			2'b11: do_bin = 2'b01;
			2'b01: do_bin = 2'b10;
			2'b00: do_bin = 2'b11;
		endcase
	end
	else begin
		case (grey[1:0])
			2'b00: do_bin = 2'b00;
			2'b01: do_bin = 2'b01;
			2'b11: do_bin = 2'b10;
			2'b10: do_bin = 2'b11;
		endcase
	end
end
endfunction
function [AW:0] get_cnt;
input [AW:0] wr_ptr, rd_ptr;
begin
	if (wr_ptr >= rd_ptr) begin
		get_cnt = (wr_ptr - rd_ptr);	
	end
	else begin
		get_cnt = DP*2 - (rd_ptr - wr_ptr);
	end
end
endfunction
// synopsys translate_off
always @(posedge wr_clk) begin
   if (wr_en && wr_full) begin
      $display($time, "%m Error! afifo overflow!");
      $stop;
   end
end
always @(posedge rd_clk) begin
   if (rd_en && rd_empty) begin
      $display($time, "%m error! afifo underflow!");
      $stop;
   end
end
// synopsys translate_on
endmodule
module ahb_matrix_1_6_sub_dec(
  hclk,
  hresetn,
  load_cmd,
  m_haddr,
  m_hburst,
  m_hprot,
  m_hrdata,
  m_hready,
  m_hresp,
  m_hsize,
  m_htrans,
  m_hwdata,
  m_hwrite,
  m_resp_vld,
  pmu_matrix_clkdiv_bypass,
  s0_haddr,
  s0_hburst,
  s0_hprot,
  s0_hrdata,
  s0_hready,
  s0_hresp,
  s0_hselx,
  s0_hsize,
  s0_htrans,
  s0_hwdata,
  s0_hwrite,
  s1_haddr,
  s1_hburst,
  s1_hprot,
  s1_hrdata,
  s1_hready,
  s1_hresp,
  s1_hselx,
  s1_hsize,
  s1_htrans,
  s1_hwdata,
  s1_hwrite,
  s2_haddr,
  s2_hburst,
  s2_hprot,
  s2_hrdata,
  s2_hready,
  s2_hresp,
  s2_hselx,
  s2_hsize,
  s2_htrans,
  s2_hwdata,
  s2_hwrite,
  s3_haddr,
  s3_hburst,
  s3_hprot,
  s3_hrdata,
  s3_hready,
  s3_hresp,
  s3_hselx,
  s3_hsize,
  s3_htrans,
  s3_hwdata,
  s3_hwrite,
  s4_haddr,
  s4_hburst,
  s4_hprot,
  s4_hrdata,
  s4_hready,
  s4_hresp,
  s4_hselx,
  s4_hsize,
  s4_htrans,
  s4_hwdata,
  s4_hwrite,
  s5_haddr,
  s5_hburst,
  s5_hprot,
  s5_hrdata,
  s5_hready,
  s5_hresp,
  s5_hselx,
  s5_hsize,
  s5_htrans,
  s5_hwdata,
  s5_hwrite,
  wfifo_rd_empty
);
input           hclk;                    
input           hresetn;                 
input   [31:0]  m_haddr;                 
input   [2 :0]  m_hburst;                
input   [3 :0]  m_hprot;                 
input   [2 :0]  m_hsize;                 
input   [1 :0]  m_htrans;                
input   [31:0]  m_hwdata;                
input           m_hwrite;                
input           pmu_matrix_clkdiv_bypass; 
input   [31:0]  s0_hrdata;               
input           s0_hready;               
input   [1 :0]  s0_hresp;                
input   [31:0]  s1_hrdata;               
input           s1_hready;               
input   [1 :0]  s1_hresp;                
input   [31:0]  s2_hrdata;               
input           s2_hready;               
input   [1 :0]  s2_hresp;                
input   [31:0]  s3_hrdata;               
input           s3_hready;               
input   [1 :0]  s3_hresp;                
input   [31:0]  s4_hrdata;               
input           s4_hready;               
input   [1 :0]  s4_hresp;                
input   [31:0]  s5_hrdata;               
input           s5_hready;               
input   [1 :0]  s5_hresp;                
input           wfifo_rd_empty;          
output          load_cmd;                
output  [31:0]  m_hrdata;                
output          m_hready;                
output  [1 :0]  m_hresp;                 
output          m_resp_vld;              
output  [31:0]  s0_haddr;                
output  [2 :0]  s0_hburst;               
output  [3 :0]  s0_hprot;                
output          s0_hselx;                
output  [2 :0]  s0_hsize;                
output  [1 :0]  s0_htrans;               
output  [31:0]  s0_hwdata;               
output          s0_hwrite;               
output  [31:0]  s1_haddr;                
output  [2 :0]  s1_hburst;               
output  [3 :0]  s1_hprot;                
output          s1_hselx;                
output  [2 :0]  s1_hsize;                
output  [1 :0]  s1_htrans;               
output  [31:0]  s1_hwdata;               
output          s1_hwrite;               
output  [31:0]  s2_haddr;                
output  [2 :0]  s2_hburst;               
output  [3 :0]  s2_hprot;                
output          s2_hselx;                
output  [2 :0]  s2_hsize;                
output  [1 :0]  s2_htrans;               
output  [31:0]  s2_hwdata;               
output          s2_hwrite;               
output  [31:0]  s3_haddr;                
output  [2 :0]  s3_hburst;               
output  [3 :0]  s3_hprot;                
output          s3_hselx;                
output  [2 :0]  s3_hsize;                
output  [1 :0]  s3_htrans;               
output  [31:0]  s3_hwdata;               
output          s3_hwrite;               
output  [31:0]  s4_haddr;                
output  [2 :0]  s4_hburst;               
output  [3 :0]  s4_hprot;                
output          s4_hselx;                
output  [2 :0]  s4_hsize;                
output  [1 :0]  s4_htrans;               
output  [31:0]  s4_hwdata;               
output          s4_hwrite;               
output  [31:0]  s5_haddr;                
output  [2 :0]  s5_hburst;               
output  [3 :0]  s5_hprot;                
output          s5_hselx;                
output  [2 :0]  s5_hsize;                
output  [1 :0]  s5_htrans;               
output  [31:0]  s5_hwdata;               
output          s5_hwrite;               
reg             clr_cmd;                 
reg             latch_cmd;               
reg             load_cmd;                
reg     [42:0]  m_ctrl_bus_d;            
reg     [12:0]  m_cur_st;                
reg             m_hready;                
reg     [31:0]  m_hwdata_d;              
reg     [12:0]  m_nxt_st;                
reg             m_resp_vld;              
reg             s0_cur_cmd;              
reg             s0_last_cmd;             
reg             s1_cur_cmd;              
reg             s1_last_cmd;             
reg             s2_cur_cmd;              
reg             s2_last_cmd;             
reg             s3_cur_cmd;              
reg             s3_last_cmd;             
reg             s4_cur_cmd;              
reg             s4_last_cmd;             
reg             s5_cur_cmd;              
reg             s5_last_cmd;             
wire            bypass_mode;             
wire            hclk;                    
wire            hresetn;                 
wire    [42:0]  m_ctrl_bus;              
wire    [31:0]  m_haddr;                 
wire    [2 :0]  m_hburst;                
wire    [3 :0]  m_hprot;                 
wire    [31:0]  m_hrdata;                
wire    [1 :0]  m_hresp;                 
wire    [2 :0]  m_hsize;                 
wire    [1 :0]  m_htrans;                
wire    [31:0]  m_hwdata;                
wire            m_hwrite;                
wire            pmu_matrix_clkdiv_bypass; 
wire    [31:0]  s0_haddr;                
wire    [2 :0]  s0_hburst;               
wire    [3 :0]  s0_hprot;                
wire    [31:0]  s0_hrdata;               
wire            s0_hready;               
wire    [1 :0]  s0_hresp;                
wire            s0_hselx;                
wire    [2 :0]  s0_hsize;                
wire    [1 :0]  s0_htrans;               
wire    [31:0]  s0_hwdata;               
wire            s0_hwrite;               
wire            s0_sel;                  
wire    [31:0]  s1_haddr;                
wire    [2 :0]  s1_hburst;               
wire    [3 :0]  s1_hprot;                
wire    [31:0]  s1_hrdata;               
wire            s1_hready;               
wire    [1 :0]  s1_hresp;                
wire            s1_hselx;                
wire    [2 :0]  s1_hsize;                
wire    [1 :0]  s1_htrans;               
wire    [31:0]  s1_hwdata;               
wire            s1_hwrite;               
wire            s1_sel;                  
wire    [31:0]  s2_haddr;                
wire    [2 :0]  s2_hburst;               
wire    [3 :0]  s2_hprot;                
wire    [31:0]  s2_hrdata;               
wire            s2_hready;               
wire    [1 :0]  s2_hresp;                
wire            s2_hselx;                
wire    [2 :0]  s2_hsize;                
wire    [1 :0]  s2_htrans;               
wire    [31:0]  s2_hwdata;               
wire            s2_hwrite;               
wire            s2_sel;                  
wire    [31:0]  s3_haddr;                
wire    [2 :0]  s3_hburst;               
wire    [3 :0]  s3_hprot;                
wire    [31:0]  s3_hrdata;               
wire            s3_hready;               
wire    [1 :0]  s3_hresp;                
wire            s3_hselx;                
wire    [2 :0]  s3_hsize;                
wire    [1 :0]  s3_htrans;               
wire    [31:0]  s3_hwdata;               
wire            s3_hwrite;               
wire            s3_sel;                  
wire    [31:0]  s4_haddr;                
wire    [2 :0]  s4_hburst;               
wire    [3 :0]  s4_hprot;                
wire    [31:0]  s4_hrdata;               
wire            s4_hready;               
wire    [1 :0]  s4_hresp;                
wire            s4_hselx;                
wire    [2 :0]  s4_hsize;                
wire    [1 :0]  s4_htrans;               
wire    [31:0]  s4_hwdata;               
wire            s4_hwrite;               
wire            s4_sel;                  
wire    [31:0]  s5_haddr;                
wire    [2 :0]  s5_hburst;               
wire    [3 :0]  s5_hprot;                
wire    [31:0]  s5_hrdata;               
wire            s5_hready;               
wire    [1 :0]  s5_hresp;                
wire            s5_hselx;                
wire    [2 :0]  s5_hsize;                
wire    [1 :0]  s5_htrans;               
wire    [31:0]  s5_hwdata;               
wire            s5_hwrite;               
wire            s5_sel;                  
wire            wfifo_rd_empty;          
parameter BUS_WIDTH = 43;
parameter S_IDLE    = 13'b0000000000001;
parameter S_S0_CMD  = 13'b0000000000010;
parameter S_S0_DATA = 13'b0000000000100;
parameter S_S1_CMD  = 13'b0000000001000;
parameter S_S1_DATA = 13'b0000000010000;
parameter S_S2_CMD  = 13'b0000000100000;
parameter S_S2_DATA = 13'b0000001000000;
parameter S_S3_CMD  = 13'b0000010000000;
parameter S_S3_DATA = 13'b0000100000000;
parameter S_S4_CMD  = 13'b0001000000000;
parameter S_S4_DATA = 13'b0010000000000;
parameter S_S5_CMD  = 13'b0100000000000;
parameter S_S5_DATA = 13'b1000000000000;
assign s0_sel =( m_haddr[31:0] >= 32'h40200000) & (m_haddr[31:0] <= 32'h40200fff) & (m_htrans[1]);
assign s1_sel =( m_haddr[31:0] >= 32'h40300000) & (m_haddr[31:0] <= 32'h403fffff) & (m_htrans[1]);
assign s2_sel =( m_haddr[31:0] >= 32'h50000000) & (m_haddr[31:0] <= 32'h5004ffff) & (m_htrans[1]);
assign s3_sel =( m_haddr[31:0] >= 32'h60000000) & (m_haddr[31:0] <= 32'h6004ffff) & (m_htrans[1]);
assign s4_sel =( m_haddr[31:0] >= 32'h70000000) & (m_haddr[31:0] <= 32'h77ffffff) & (m_htrans[1]);
assign s5_sel =( m_haddr[31:0] >= 32'h78000000) & (m_haddr[31:0] <= 32'h7fffffff) & (m_htrans[1]);
assign bypass_mode = pmu_matrix_clkdiv_bypass;
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
       m_cur_st[12:0] <= S_IDLE;
    else
       m_cur_st[12:0] <= m_nxt_st[12:0];
  end
always @ (*)
begin
case(m_cur_st[12:0])
  S_IDLE:begin
       load_cmd = bypass_mode ? 1'b0 : ~wfifo_rd_empty;
       clr_cmd = 1'b0;
       m_resp_vld = 1'b0;
       latch_cmd = 1'b0;
       s0_cur_cmd = 1'b0;
       s0_last_cmd = 1'b0;
       s1_cur_cmd = 1'b0;
       s1_last_cmd = 1'b0;
       s2_cur_cmd = 1'b0;
       s2_last_cmd = 1'b0;
       s3_cur_cmd = 1'b0;
       s3_last_cmd = 1'b0;
       s4_cur_cmd = 1'b0;
       s4_last_cmd = 1'b0;
       s5_cur_cmd = 1'b0;
       s5_last_cmd = 1'b0;
       case(1'b1)
         s0_sel: begin 
                   m_nxt_st[12:0] = bypass_mode ? (s0_hready ? S_S0_DATA : S_S0_CMD) : S_S0_CMD;
                   s0_cur_cmd = bypass_mode ? (s0_hready ? 1'b1 : 1'b0) : 1'b0;
                   latch_cmd = bypass_mode ? (s0_hready ? 1'b0 : 1'b1) : 1'b0;
         end
         s1_sel: begin 
                   m_nxt_st[12:0] = bypass_mode ? (s1_hready ? S_S1_DATA : S_S1_CMD) : S_S1_CMD;
                   s1_cur_cmd = bypass_mode ? (s1_hready ? 1'b1 : 1'b0) : 1'b0;
                   latch_cmd = bypass_mode ? (s1_hready ? 1'b0 : 1'b1) : 1'b0;
         end
         s2_sel: begin 
                   m_nxt_st[12:0] = bypass_mode ? (s2_hready ? S_S2_DATA : S_S2_CMD) : S_S2_CMD;
                   s2_cur_cmd = bypass_mode ? (s2_hready ? 1'b1 : 1'b0) : 1'b0;
                   latch_cmd = bypass_mode ? (s2_hready ? 1'b0 : 1'b1) : 1'b0;
         end
         s3_sel: begin 
                   m_nxt_st[12:0] = bypass_mode ? (s3_hready ? S_S3_DATA : S_S3_CMD) : S_S3_CMD;
                   s3_cur_cmd = bypass_mode ? (s3_hready ? 1'b1 : 1'b0) : 1'b0;
                   latch_cmd = bypass_mode ? (s3_hready ? 1'b0 : 1'b1) : 1'b0;
         end
         s4_sel: begin 
                   m_nxt_st[12:0] = bypass_mode ? (s4_hready ? S_S4_DATA : S_S4_CMD) : S_S4_CMD;
                   s4_cur_cmd = bypass_mode ? (s4_hready ? 1'b1 : 1'b0) : 1'b0;
                   latch_cmd = bypass_mode ? (s4_hready ? 1'b0 : 1'b1) : 1'b0;
         end
         s5_sel: begin 
                   m_nxt_st[12:0] = bypass_mode ? (s5_hready ? S_S5_DATA : S_S5_CMD) : S_S5_CMD;
                   s5_cur_cmd = bypass_mode ? (s5_hready ? 1'b1 : 1'b0) : 1'b0;
                   latch_cmd = bypass_mode ? (s5_hready ? 1'b0 : 1'b1) : 1'b0;
         end
         default: m_nxt_st[12:0] = S_IDLE;
       endcase
  end
  S_S0_CMD:begin
     load_cmd = 1'b0;
     clr_cmd = s0_hready ? 1'b1 : 1'b0;
     s0_cur_cmd = 1'b0;
     s0_last_cmd = 1'b1;
     s1_cur_cmd = 1'b0;
     s1_last_cmd = 1'b0;
     s2_cur_cmd = 1'b0;
     s2_last_cmd = 1'b0;
     s3_cur_cmd = 1'b0;
     s3_last_cmd = 1'b0;
     s4_cur_cmd = 1'b0;
     s4_last_cmd = 1'b0;
     s5_cur_cmd = 1'b0;
     s5_last_cmd = 1'b0;
     latch_cmd = 1'b0;
     m_resp_vld = 1'b0;
     m_nxt_st[12:0] = s0_hready ? S_S0_DATA : S_S0_CMD;
  end
  S_S0_DATA:begin
     load_cmd = 1'b0;
     clr_cmd = 1'b0;
     s0_cur_cmd = 1'b0;
     s0_last_cmd = 1'b0;
     s1_cur_cmd = 1'b0;
     s1_last_cmd = 1'b0;
     s2_cur_cmd = 1'b0;
     s2_last_cmd = 1'b0;
     s3_cur_cmd = 1'b0;
     s3_last_cmd = 1'b0;
     s4_cur_cmd = 1'b0;
     s4_last_cmd = 1'b0;
     s5_cur_cmd = 1'b0;
     s5_last_cmd = 1'b0;
     latch_cmd = 1'b0;
     m_resp_vld = 1'b0;
     if(s0_hready) begin
       load_cmd = bypass_mode ? 1'b0 : ~wfifo_rd_empty;
       m_resp_vld = 1'b1;
       case(1'b1)
         s0_sel: begin 
                   m_nxt_st[12:0] = s0_hready ? S_S0_DATA : S_S0_CMD;
                   latch_cmd = s0_hready ? 1'b0 : 1'b1;
                   s0_cur_cmd = s0_hready  ? 1'b1 : 1'b0;
         end
         s1_sel: begin 
                   m_nxt_st[12:0] = s1_hready ? S_S1_DATA : S_S1_CMD;
                   latch_cmd = s1_hready ? 1'b0 : 1'b1;
                   s1_cur_cmd = s1_hready  ? 1'b1 : 1'b0;
         end
         s2_sel: begin 
                   m_nxt_st[12:0] = s2_hready ? S_S2_DATA : S_S2_CMD;
                   latch_cmd = s2_hready ? 1'b0 : 1'b1;
                   s2_cur_cmd = s2_hready  ? 1'b1 : 1'b0;
         end
         s3_sel: begin 
                   m_nxt_st[12:0] = s3_hready ? S_S3_DATA : S_S3_CMD;
                   latch_cmd = s3_hready ? 1'b0 : 1'b1;
                   s3_cur_cmd = s3_hready  ? 1'b1 : 1'b0;
         end
         s4_sel: begin 
                   m_nxt_st[12:0] = s4_hready ? S_S4_DATA : S_S4_CMD;
                   latch_cmd = s4_hready ? 1'b0 : 1'b1;
                   s4_cur_cmd = s4_hready  ? 1'b1 : 1'b0;
         end
         s5_sel: begin 
                   m_nxt_st[12:0] = s5_hready ? S_S5_DATA : S_S5_CMD;
                   latch_cmd = s5_hready ? 1'b0 : 1'b1;
                   s5_cur_cmd = s5_hready  ? 1'b1 : 1'b0;
         end
         default: m_nxt_st[12:0] = S_IDLE;
       endcase
     end
     else begin
       m_nxt_st[12:0] = S_S0_DATA;
     end
  end
  S_S1_CMD:begin
     load_cmd = 1'b0;
     clr_cmd = s1_hready ? 1'b1 : 1'b0;
     s0_cur_cmd = 1'b0;
     s0_last_cmd = 1'b0;
     s1_cur_cmd = 1'b0;
     s1_last_cmd = 1'b1;
     s2_cur_cmd = 1'b0;
     s2_last_cmd = 1'b0;
     s3_cur_cmd = 1'b0;
     s3_last_cmd = 1'b0;
     s4_cur_cmd = 1'b0;
     s4_last_cmd = 1'b0;
     s5_cur_cmd = 1'b0;
     s5_last_cmd = 1'b0;
     latch_cmd = 1'b0;
     m_resp_vld = 1'b0;
     m_nxt_st[12:0] = s1_hready ? S_S1_DATA : S_S1_CMD;
  end
  S_S1_DATA:begin
     load_cmd = 1'b0;
     clr_cmd = 1'b0;
     s0_cur_cmd = 1'b0;
     s0_last_cmd = 1'b0;
     s1_cur_cmd = 1'b0;
     s1_last_cmd = 1'b0;
     s2_cur_cmd = 1'b0;
     s2_last_cmd = 1'b0;
     s3_cur_cmd = 1'b0;
     s3_last_cmd = 1'b0;
     s4_cur_cmd = 1'b0;
     s4_last_cmd = 1'b0;
     s5_cur_cmd = 1'b0;
     s5_last_cmd = 1'b0;
     latch_cmd = 1'b0;
     m_resp_vld = 1'b0;
     if(s1_hready) begin
       load_cmd = bypass_mode ? 1'b0 : ~wfifo_rd_empty;
       m_resp_vld = 1'b1;
       case(1'b1)
         s0_sel: begin 
                   m_nxt_st[12:0] = s0_hready ? S_S0_DATA : S_S0_CMD;
                   latch_cmd = s0_hready ? 1'b0 : 1'b1;
                   s0_cur_cmd = s0_hready  ? 1'b1 : 1'b0;
         end
         s1_sel: begin 
                   m_nxt_st[12:0] = s1_hready ? S_S1_DATA : S_S1_CMD;
                   latch_cmd = s1_hready ? 1'b0 : 1'b1;
                   s1_cur_cmd = s1_hready  ? 1'b1 : 1'b0;
         end
         s2_sel: begin 
                   m_nxt_st[12:0] = s2_hready ? S_S2_DATA : S_S2_CMD;
                   latch_cmd = s2_hready ? 1'b0 : 1'b1;
                   s2_cur_cmd = s2_hready  ? 1'b1 : 1'b0;
         end
         s3_sel: begin 
                   m_nxt_st[12:0] = s3_hready ? S_S3_DATA : S_S3_CMD;
                   latch_cmd = s3_hready ? 1'b0 : 1'b1;
                   s3_cur_cmd = s3_hready  ? 1'b1 : 1'b0;
         end
         s4_sel: begin 
                   m_nxt_st[12:0] = s4_hready ? S_S4_DATA : S_S4_CMD;
                   latch_cmd = s4_hready ? 1'b0 : 1'b1;
                   s4_cur_cmd = s4_hready  ? 1'b1 : 1'b0;
         end
         s5_sel: begin 
                   m_nxt_st[12:0] = s5_hready ? S_S5_DATA : S_S5_CMD;
                   latch_cmd = s5_hready ? 1'b0 : 1'b1;
                   s5_cur_cmd = s5_hready  ? 1'b1 : 1'b0;
         end
         default: m_nxt_st[12:0] = S_IDLE;
       endcase
     end
     else begin
       m_nxt_st[12:0] = S_S1_DATA;
     end
  end
  S_S2_CMD:begin
     load_cmd = 1'b0;
     clr_cmd = s2_hready ? 1'b1 : 1'b0;
     s0_cur_cmd = 1'b0;
     s0_last_cmd = 1'b0;
     s1_cur_cmd = 1'b0;
     s1_last_cmd = 1'b0;
     s2_cur_cmd = 1'b0;
     s2_last_cmd = 1'b1;
     s3_cur_cmd = 1'b0;
     s3_last_cmd = 1'b0;
     s4_cur_cmd = 1'b0;
     s4_last_cmd = 1'b0;
     s5_cur_cmd = 1'b0;
     s5_last_cmd = 1'b0;
     latch_cmd = 1'b0;
     m_resp_vld = 1'b0;
     m_nxt_st[12:0] = s2_hready ? S_S2_DATA : S_S2_CMD;
  end
  S_S2_DATA:begin
     load_cmd = 1'b0;
     clr_cmd = 1'b0;
     s0_cur_cmd = 1'b0;
     s0_last_cmd = 1'b0;
     s1_cur_cmd = 1'b0;
     s1_last_cmd = 1'b0;
     s2_cur_cmd = 1'b0;
     s2_last_cmd = 1'b0;
     s3_cur_cmd = 1'b0;
     s3_last_cmd = 1'b0;
     s4_cur_cmd = 1'b0;
     s4_last_cmd = 1'b0;
     s5_cur_cmd = 1'b0;
     s5_last_cmd = 1'b0;
     latch_cmd = 1'b0;
     m_resp_vld = 1'b0;
     if(s2_hready) begin
       load_cmd = bypass_mode ? 1'b0 : ~wfifo_rd_empty;
       m_resp_vld = 1'b1;
       case(1'b1)
         s0_sel: begin 
                   m_nxt_st[12:0] = s0_hready ? S_S0_DATA : S_S0_CMD;
                   latch_cmd = s0_hready ? 1'b0 : 1'b1;
                   s0_cur_cmd = s0_hready  ? 1'b1 : 1'b0;
         end
         s1_sel: begin 
                   m_nxt_st[12:0] = s1_hready ? S_S1_DATA : S_S1_CMD;
                   latch_cmd = s1_hready ? 1'b0 : 1'b1;
                   s1_cur_cmd = s1_hready  ? 1'b1 : 1'b0;
         end
         s2_sel: begin 
                   m_nxt_st[12:0] = s2_hready ? S_S2_DATA : S_S2_CMD;
                   latch_cmd = s2_hready ? 1'b0 : 1'b1;
                   s2_cur_cmd = s2_hready  ? 1'b1 : 1'b0;
         end
         s3_sel: begin 
                   m_nxt_st[12:0] = s3_hready ? S_S3_DATA : S_S3_CMD;
                   latch_cmd = s3_hready ? 1'b0 : 1'b1;
                   s3_cur_cmd = s3_hready  ? 1'b1 : 1'b0;
         end
         s4_sel: begin 
                   m_nxt_st[12:0] = s4_hready ? S_S4_DATA : S_S4_CMD;
                   latch_cmd = s4_hready ? 1'b0 : 1'b1;
                   s4_cur_cmd = s4_hready  ? 1'b1 : 1'b0;
         end
         s5_sel: begin 
                   m_nxt_st[12:0] = s5_hready ? S_S5_DATA : S_S5_CMD;
                   latch_cmd = s5_hready ? 1'b0 : 1'b1;
                   s5_cur_cmd = s5_hready  ? 1'b1 : 1'b0;
         end
         default: m_nxt_st[12:0] = S_IDLE;
       endcase
     end
     else begin
       m_nxt_st[12:0] = S_S2_DATA;
     end
  end
  S_S3_CMD:begin
     load_cmd = 1'b0;
     clr_cmd = s3_hready ? 1'b1 : 1'b0;
     s0_cur_cmd = 1'b0;
     s0_last_cmd = 1'b0;
     s1_cur_cmd = 1'b0;
     s1_last_cmd = 1'b0;
     s2_cur_cmd = 1'b0;
     s2_last_cmd = 1'b0;
     s3_cur_cmd = 1'b0;
     s3_last_cmd = 1'b1;
     s4_cur_cmd = 1'b0;
     s4_last_cmd = 1'b0;
     s5_cur_cmd = 1'b0;
     s5_last_cmd = 1'b0;
     latch_cmd = 1'b0;
     m_resp_vld = 1'b0;
     m_nxt_st[12:0] = s3_hready ? S_S3_DATA : S_S3_CMD;
  end
  S_S3_DATA:begin
     load_cmd = 1'b0;
     clr_cmd = 1'b0;
     s0_cur_cmd = 1'b0;
     s0_last_cmd = 1'b0;
     s1_cur_cmd = 1'b0;
     s1_last_cmd = 1'b0;
     s2_cur_cmd = 1'b0;
     s2_last_cmd = 1'b0;
     s3_cur_cmd = 1'b0;
     s3_last_cmd = 1'b0;
     s4_cur_cmd = 1'b0;
     s4_last_cmd = 1'b0;
     s5_cur_cmd = 1'b0;
     s5_last_cmd = 1'b0;
     latch_cmd = 1'b0;
     m_resp_vld = 1'b0;
     if(s3_hready) begin
       load_cmd = bypass_mode ? 1'b0 : ~wfifo_rd_empty;
       m_resp_vld = 1'b1;
       case(1'b1)
         s0_sel: begin 
                   m_nxt_st[12:0] = s0_hready ? S_S0_DATA : S_S0_CMD;
                   latch_cmd = s0_hready ? 1'b0 : 1'b1;
                   s0_cur_cmd = s0_hready  ? 1'b1 : 1'b0;
         end
         s1_sel: begin 
                   m_nxt_st[12:0] = s1_hready ? S_S1_DATA : S_S1_CMD;
                   latch_cmd = s1_hready ? 1'b0 : 1'b1;
                   s1_cur_cmd = s1_hready  ? 1'b1 : 1'b0;
         end
         s2_sel: begin 
                   m_nxt_st[12:0] = s2_hready ? S_S2_DATA : S_S2_CMD;
                   latch_cmd = s2_hready ? 1'b0 : 1'b1;
                   s2_cur_cmd = s2_hready  ? 1'b1 : 1'b0;
         end
         s3_sel: begin 
                   m_nxt_st[12:0] = s3_hready ? S_S3_DATA : S_S3_CMD;
                   latch_cmd = s3_hready ? 1'b0 : 1'b1;
                   s3_cur_cmd = s3_hready  ? 1'b1 : 1'b0;
         end
         s4_sel: begin 
                   m_nxt_st[12:0] = s4_hready ? S_S4_DATA : S_S4_CMD;
                   latch_cmd = s4_hready ? 1'b0 : 1'b1;
                   s4_cur_cmd = s4_hready  ? 1'b1 : 1'b0;
         end
         s5_sel: begin 
                   m_nxt_st[12:0] = s5_hready ? S_S5_DATA : S_S5_CMD;
                   latch_cmd = s5_hready ? 1'b0 : 1'b1;
                   s5_cur_cmd = s5_hready  ? 1'b1 : 1'b0;
         end
         default: m_nxt_st[12:0] = S_IDLE;
       endcase
     end
     else begin
       m_nxt_st[12:0] = S_S3_DATA;
     end
  end
  S_S4_CMD:begin
     load_cmd = 1'b0;
     clr_cmd = s4_hready ? 1'b1 : 1'b0;
     s0_cur_cmd = 1'b0;
     s0_last_cmd = 1'b0;
     s1_cur_cmd = 1'b0;
     s1_last_cmd = 1'b0;
     s2_cur_cmd = 1'b0;
     s2_last_cmd = 1'b0;
     s3_cur_cmd = 1'b0;
     s3_last_cmd = 1'b0;
     s4_cur_cmd = 1'b0;
     s4_last_cmd = 1'b1;
     s5_cur_cmd = 1'b0;
     s5_last_cmd = 1'b0;
     latch_cmd = 1'b0;
     m_resp_vld = 1'b0;
     m_nxt_st[12:0] = s4_hready ? S_S4_DATA : S_S4_CMD;
  end
  S_S4_DATA:begin
     load_cmd = 1'b0;
     clr_cmd = 1'b0;
     s0_cur_cmd = 1'b0;
     s0_last_cmd = 1'b0;
     s1_cur_cmd = 1'b0;
     s1_last_cmd = 1'b0;
     s2_cur_cmd = 1'b0;
     s2_last_cmd = 1'b0;
     s3_cur_cmd = 1'b0;
     s3_last_cmd = 1'b0;
     s4_cur_cmd = 1'b0;
     s4_last_cmd = 1'b0;
     s5_cur_cmd = 1'b0;
     s5_last_cmd = 1'b0;
     latch_cmd = 1'b0;
     m_resp_vld = 1'b0;
     if(s4_hready) begin
       load_cmd = bypass_mode ? 1'b0 : ~wfifo_rd_empty;
       m_resp_vld = 1'b1;
       case(1'b1)
         s0_sel: begin 
                   m_nxt_st[12:0] = s0_hready ? S_S0_DATA : S_S0_CMD;
                   latch_cmd = s0_hready ? 1'b0 : 1'b1;
                   s0_cur_cmd = s0_hready  ? 1'b1 : 1'b0;
         end
         s1_sel: begin 
                   m_nxt_st[12:0] = s1_hready ? S_S1_DATA : S_S1_CMD;
                   latch_cmd = s1_hready ? 1'b0 : 1'b1;
                   s1_cur_cmd = s1_hready  ? 1'b1 : 1'b0;
         end
         s2_sel: begin 
                   m_nxt_st[12:0] = s2_hready ? S_S2_DATA : S_S2_CMD;
                   latch_cmd = s2_hready ? 1'b0 : 1'b1;
                   s2_cur_cmd = s2_hready  ? 1'b1 : 1'b0;
         end
         s3_sel: begin 
                   m_nxt_st[12:0] = s3_hready ? S_S3_DATA : S_S3_CMD;
                   latch_cmd = s3_hready ? 1'b0 : 1'b1;
                   s3_cur_cmd = s3_hready  ? 1'b1 : 1'b0;
         end
         s4_sel: begin 
                   m_nxt_st[12:0] = s4_hready ? S_S4_DATA : S_S4_CMD;
                   latch_cmd = s4_hready ? 1'b0 : 1'b1;
                   s4_cur_cmd = s4_hready  ? 1'b1 : 1'b0;
         end
         s5_sel: begin 
                   m_nxt_st[12:0] = s5_hready ? S_S5_DATA : S_S5_CMD;
                   latch_cmd = s5_hready ? 1'b0 : 1'b1;
                   s5_cur_cmd = s5_hready  ? 1'b1 : 1'b0;
         end
         default: m_nxt_st[12:0] = S_IDLE;
       endcase
     end
     else begin
       m_nxt_st[12:0] = S_S4_DATA;
     end
  end
  S_S5_CMD:begin
     load_cmd = 1'b0;
     clr_cmd = s5_hready ? 1'b1 : 1'b0;
     s0_cur_cmd = 1'b0;
     s0_last_cmd = 1'b0;
     s1_cur_cmd = 1'b0;
     s1_last_cmd = 1'b0;
     s2_cur_cmd = 1'b0;
     s2_last_cmd = 1'b0;
     s3_cur_cmd = 1'b0;
     s3_last_cmd = 1'b0;
     s4_cur_cmd = 1'b0;
     s4_last_cmd = 1'b0;
     s5_cur_cmd = 1'b0;
     s5_last_cmd = 1'b1;
     latch_cmd = 1'b0;
     m_resp_vld = 1'b0;
     m_nxt_st[12:0] = s5_hready ? S_S5_DATA : S_S5_CMD;
  end
  S_S5_DATA:begin
     load_cmd = 1'b0;
     clr_cmd = 1'b0;
     s0_cur_cmd = 1'b0;
     s0_last_cmd = 1'b0;
     s1_cur_cmd = 1'b0;
     s1_last_cmd = 1'b0;
     s2_cur_cmd = 1'b0;
     s2_last_cmd = 1'b0;
     s3_cur_cmd = 1'b0;
     s3_last_cmd = 1'b0;
     s4_cur_cmd = 1'b0;
     s4_last_cmd = 1'b0;
     s5_cur_cmd = 1'b0;
     s5_last_cmd = 1'b0;
     latch_cmd = 1'b0;
     m_resp_vld = 1'b0;
     if(s5_hready) begin
       load_cmd = bypass_mode ? 1'b0 : ~wfifo_rd_empty;
       m_resp_vld = 1'b1;
       case(1'b1)
         s0_sel: begin 
                   m_nxt_st[12:0] = s0_hready ? S_S0_DATA : S_S0_CMD;
                   latch_cmd = s0_hready ? 1'b0 : 1'b1;
                   s0_cur_cmd = s0_hready  ? 1'b1 : 1'b0;
         end
         s1_sel: begin 
                   m_nxt_st[12:0] = s1_hready ? S_S1_DATA : S_S1_CMD;
                   latch_cmd = s1_hready ? 1'b0 : 1'b1;
                   s1_cur_cmd = s1_hready  ? 1'b1 : 1'b0;
         end
         s2_sel: begin 
                   m_nxt_st[12:0] = s2_hready ? S_S2_DATA : S_S2_CMD;
                   latch_cmd = s2_hready ? 1'b0 : 1'b1;
                   s2_cur_cmd = s2_hready  ? 1'b1 : 1'b0;
         end
         s3_sel: begin 
                   m_nxt_st[12:0] = s3_hready ? S_S3_DATA : S_S3_CMD;
                   latch_cmd = s3_hready ? 1'b0 : 1'b1;
                   s3_cur_cmd = s3_hready  ? 1'b1 : 1'b0;
         end
         s4_sel: begin 
                   m_nxt_st[12:0] = s4_hready ? S_S4_DATA : S_S4_CMD;
                   latch_cmd = s4_hready ? 1'b0 : 1'b1;
                   s4_cur_cmd = s4_hready  ? 1'b1 : 1'b0;
         end
         s5_sel: begin 
                   m_nxt_st[12:0] = s5_hready ? S_S5_DATA : S_S5_CMD;
                   latch_cmd = s5_hready ? 1'b0 : 1'b1;
                   s5_cur_cmd = s5_hready  ? 1'b1 : 1'b0;
         end
         default: m_nxt_st[12:0] = S_IDLE;
       endcase
     end
     else begin
       m_nxt_st[12:0] = S_S5_DATA;
     end
  end
  default: begin
             m_nxt_st[12:0] = S_IDLE;
             load_cmd = bypass_mode ? 1'b0 : ~wfifo_rd_empty;
             clr_cmd = 1'b0;
             m_resp_vld = 1'b0;
             latch_cmd = 1'b0;
             s0_cur_cmd = 1'b0;
             s0_last_cmd = 1'b0;
             s1_cur_cmd = 1'b0;
             s1_last_cmd = 1'b0;
             s2_cur_cmd = 1'b0;
             s2_last_cmd = 1'b0;
             s3_cur_cmd = 1'b0;
             s3_last_cmd = 1'b0;
             s4_cur_cmd = 1'b0;
             s4_last_cmd = 1'b0;
             s5_cur_cmd = 1'b0;
             s5_last_cmd = 1'b0;
  end
endcase
end
assign m_ctrl_bus[BUS_WIDTH-1:0] = {m_haddr[32-1:0],m_hsize[2:0],m_hburst[2:0],m_hprot[3:0],m_hwrite};
assign {s0_haddr[32-1:0],s0_hsize[2:0],s0_hburst[2:0],s0_hprot[3:0],s0_hwrite} = s0_cur_cmd ? m_ctrl_bus[BUS_WIDTH-1:0] : m_ctrl_bus_d[BUS_WIDTH-1:0];
assign s0_htrans[1:0] = (s0_cur_cmd | s0_last_cmd) ? 2'b10 : 2'b00;
assign {s1_haddr[32-1:0],s1_hsize[2:0],s1_hburst[2:0],s1_hprot[3:0],s1_hwrite} = s1_cur_cmd ? m_ctrl_bus[BUS_WIDTH-1:0] : m_ctrl_bus_d[BUS_WIDTH-1:0];
assign s1_htrans[1:0] = (s1_cur_cmd | s1_last_cmd) ? 2'b10 : 2'b00;
assign {s2_haddr[32-1:0],s2_hsize[2:0],s2_hburst[2:0],s2_hprot[3:0],s2_hwrite} = s2_cur_cmd ? m_ctrl_bus[BUS_WIDTH-1:0] : m_ctrl_bus_d[BUS_WIDTH-1:0];
assign s2_htrans[1:0] = (s2_cur_cmd | s2_last_cmd) ? 2'b10 : 2'b00;
assign {s3_haddr[32-1:0],s3_hsize[2:0],s3_hburst[2:0],s3_hprot[3:0],s3_hwrite} = s3_cur_cmd ? m_ctrl_bus[BUS_WIDTH-1:0] : m_ctrl_bus_d[BUS_WIDTH-1:0];
assign s3_htrans[1:0] = (s3_cur_cmd | s3_last_cmd) ? 2'b10 : 2'b00;
assign {s4_haddr[32-1:0],s4_hsize[2:0],s4_hburst[2:0],s4_hprot[3:0],s4_hwrite} = s4_cur_cmd ? m_ctrl_bus[BUS_WIDTH-1:0] : m_ctrl_bus_d[BUS_WIDTH-1:0];
assign s4_htrans[1:0] = (s4_cur_cmd | s4_last_cmd) ? 2'b10 : 2'b00;
assign {s5_haddr[32-1:0],s5_hsize[2:0],s5_hburst[2:0],s5_hprot[3:0],s5_hwrite} = s5_cur_cmd ? m_ctrl_bus[BUS_WIDTH-1:0] : m_ctrl_bus_d[BUS_WIDTH-1:0];
assign s5_htrans[1:0] = (s5_cur_cmd | s5_last_cmd) ? 2'b10 : 2'b00;
always @ (posedge hclk or negedge hresetn)
    begin
      if(!hresetn) begin
        m_ctrl_bus_d[BUS_WIDTH-1:0] <= 0;
        m_hwdata_d[32-1:0] <= 0;
      end
      else if (load_cmd | latch_cmd) begin
        m_ctrl_bus_d[BUS_WIDTH-1:0] <= m_ctrl_bus[BUS_WIDTH-1:0];
        m_hwdata_d[32-1:0] <= m_hwdata[32-1:0];
      end
      else if (clr_cmd) begin
        m_ctrl_bus_d[BUS_WIDTH-1:0] <= 0;
        m_hwdata_d[32-1:0] <= m_hwdata_d[32-1:0];
      end
    end
assign s0_hwdata[32-1:0] = m_cur_st[2] ? (bypass_mode ? m_hwdata[32-1:0] : m_hwdata_d[32-1:0] ): 0;
assign s1_hwdata[32-1:0] = m_cur_st[4] ? (bypass_mode ? m_hwdata[32-1:0] : m_hwdata_d[32-1:0] ): 0;
assign s2_hwdata[32-1:0] = m_cur_st[6] ? (bypass_mode ? m_hwdata[32-1:0] : m_hwdata_d[32-1:0] ): 0;
assign s3_hwdata[32-1:0] = m_cur_st[8] ? (bypass_mode ? m_hwdata[32-1:0] : m_hwdata_d[32-1:0] ): 0;
assign s4_hwdata[32-1:0] = m_cur_st[10] ? (bypass_mode ? m_hwdata[32-1:0] : m_hwdata_d[32-1:0] ): 0;
assign s5_hwdata[32-1:0] = m_cur_st[12] ? (bypass_mode ? m_hwdata[32-1:0] : m_hwdata_d[32-1:0] ): 0;
assign m_hrdata[32-1:0] = 
                           (s0_hrdata[32-1:0] & {32{m_cur_st[2]}}) |
                           (s1_hrdata[32-1:0] & {32{m_cur_st[4]}}) |
                           (s2_hrdata[32-1:0] & {32{m_cur_st[6]}}) |
                           (s3_hrdata[32-1:0] & {32{m_cur_st[8]}}) |
                           (s4_hrdata[32-1:0] & {32{m_cur_st[10]}}) |
                           (s5_hrdata[32-1:0] & {32{m_cur_st[12]}});
assign m_hresp[1:0] = 
                       (s0_hresp[1:0] & {2{m_cur_st[2]}}) |
                       (s1_hresp[1:0] & {2{m_cur_st[4]}}) |
                       (s2_hresp[1:0] & {2{m_cur_st[6]}}) |
                       (s3_hresp[1:0] & {2{m_cur_st[8]}}) |
                       (s4_hresp[1:0] & {2{m_cur_st[10]}}) |
                       (s5_hresp[1:0] & {2{m_cur_st[12]}});
always @( s4_hready
       or s2_hready
       or m_cur_st[12:0]
       or s1_hready
       or s3_hready
       or s5_hready
       or s0_hready)
begin
case(m_cur_st[12:0])
   S_IDLE : m_hready = 1'b1;
   S_S0_CMD: m_hready = 1'b0;
   S_S1_CMD: m_hready = 1'b0;
   S_S2_CMD: m_hready = 1'b0;
   S_S3_CMD: m_hready = 1'b0;
   S_S4_CMD: m_hready = 1'b0;
   S_S5_CMD: m_hready = 1'b0;
   S_S0_DATA: m_hready = s0_hready;
   S_S1_DATA: m_hready = s1_hready;
   S_S2_DATA: m_hready = s2_hready;
   S_S3_DATA: m_hready = s3_hready;
   S_S4_DATA: m_hready = s4_hready;
   S_S5_DATA: m_hready = s5_hready;
   default: m_hready = 1'b1;
endcase
end
assign s0_hselx = s0_cur_cmd | s0_last_cmd ;
assign s1_hselx = s1_cur_cmd | s1_last_cmd ;
assign s2_hselx = s2_cur_cmd | s2_last_cmd ;
assign s3_hselx = s3_cur_cmd | s3_last_cmd ;
assign s4_hselx = s4_cur_cmd | s4_last_cmd ;
assign s5_hselx = s5_cur_cmd | s5_last_cmd ;
endmodule
module ahb_matrix_1_6_sub(
  m_haddr,
  m_hburst,
  m_hprot,
  m_hrdata,
  m_hready,
  m_hresp,
  m_hselx,
  m_hsize,
  m_htrans,
  m_hwdata,
  m_hwrite,
  main_hclk,
  main_hresetn,
  pmu_matrix_clkdiv_bypass,
  s0_haddr,
  s0_hburst,
  s0_hprot,
  s0_hrdata,
  s0_hready,
  s0_hresp,
  s0_hselx,
  s0_hsize,
  s0_htrans,
  s0_hwdata,
  s0_hwrite,
  s1_haddr,
  s1_hburst,
  s1_hprot,
  s1_hrdata,
  s1_hready,
  s1_hresp,
  s1_hselx,
  s1_hsize,
  s1_htrans,
  s1_hwdata,
  s1_hwrite,
  s2_haddr,
  s2_hburst,
  s2_hprot,
  s2_hrdata,
  s2_hready,
  s2_hresp,
  s2_hselx,
  s2_hsize,
  s2_htrans,
  s2_hwdata,
  s2_hwrite,
  s3_haddr,
  s3_hburst,
  s3_hprot,
  s3_hrdata,
  s3_hready,
  s3_hresp,
  s3_hselx,
  s3_hsize,
  s3_htrans,
  s3_hwdata,
  s3_hwrite,
  s4_haddr,
  s4_hburst,
  s4_hprot,
  s4_hrdata,
  s4_hready,
  s4_hresp,
  s4_hselx,
  s4_hsize,
  s4_htrans,
  s4_hwdata,
  s4_hwrite,
  s5_haddr,
  s5_hburst,
  s5_hprot,
  s5_hrdata,
  s5_hready,
  s5_hresp,
  s5_hselx,
  s5_hsize,
  s5_htrans,
  s5_hwdata,
  s5_hwrite,
  sub_hclk,
  sub_hresetn
);
input   [31:0]  m_haddr;                 
input   [2 :0]  m_hburst;                
input   [3 :0]  m_hprot;                 
input           m_hselx;                 
input   [2 :0]  m_hsize;                 
input   [1 :0]  m_htrans;                
input   [31:0]  m_hwdata;                
input           m_hwrite;                
input           main_hclk;               
input           main_hresetn;            
input           pmu_matrix_clkdiv_bypass; 
input   [31:0]  s0_hrdata;               
input           s0_hready;               
input   [1 :0]  s0_hresp;                
input   [31:0]  s1_hrdata;               
input           s1_hready;               
input   [1 :0]  s1_hresp;                
input   [31:0]  s2_hrdata;               
input           s2_hready;               
input   [1 :0]  s2_hresp;                
input   [31:0]  s3_hrdata;               
input           s3_hready;               
input   [1 :0]  s3_hresp;                
input   [31:0]  s4_hrdata;               
input           s4_hready;               
input   [1 :0]  s4_hresp;                
input   [31:0]  s5_hrdata;               
input           s5_hready;               
input   [1 :0]  s5_hresp;                
input           sub_hclk;                
input           sub_hresetn;             
output  [31:0]  m_hrdata;                
output          m_hready;                
output  [1 :0]  m_hresp;                 
output  [31:0]  s0_haddr;                
output  [2 :0]  s0_hburst;               
output  [3 :0]  s0_hprot;                
output          s0_hselx;                
output  [2 :0]  s0_hsize;                
output  [1 :0]  s0_htrans;               
output  [31:0]  s0_hwdata;               
output          s0_hwrite;               
output  [31:0]  s1_haddr;                
output  [2 :0]  s1_hburst;               
output  [3 :0]  s1_hprot;                
output          s1_hselx;                
output  [2 :0]  s1_hsize;                
output  [1 :0]  s1_htrans;               
output  [31:0]  s1_hwdata;               
output          s1_hwrite;               
output  [31:0]  s2_haddr;                
output  [2 :0]  s2_hburst;               
output  [3 :0]  s2_hprot;                
output          s2_hselx;                
output  [2 :0]  s2_hsize;                
output  [1 :0]  s2_htrans;               
output  [31:0]  s2_hwdata;               
output          s2_hwrite;               
output  [31:0]  s3_haddr;                
output  [2 :0]  s3_hburst;               
output  [3 :0]  s3_hprot;                
output          s3_hselx;                
output  [2 :0]  s3_hsize;                
output  [1 :0]  s3_htrans;               
output  [31:0]  s3_hwdata;               
output          s3_hwrite;               
output  [31:0]  s4_haddr;                
output  [2 :0]  s4_hburst;               
output  [3 :0]  s4_hprot;                
output          s4_hselx;                
output  [2 :0]  s4_hsize;                
output  [1 :0]  s4_htrans;               
output  [31:0]  s4_hwdata;               
output          s4_hwrite;               
output  [31:0]  s5_haddr;                
output  [2 :0]  s5_hburst;               
output  [3 :0]  s5_hprot;                
output          s5_hselx;                
output  [2 :0]  s5_hsize;                
output  [1 :0]  s5_htrans;               
output  [31:0]  s5_hwdata;               
output          s5_hwrite;               
reg             clk_div;                 
reg     [31:0]  m_haddr_d;               
reg     [2 :0]  m_hburst_d;              
reg     [3 :0]  m_hprot_d;               
reg     [2 :0]  m_hsize_d;               
reg     [1 :0]  m_htrans_d;              
reg             m_hwrite_d;              
reg             rd_hready;               
reg             wfifo_wr_en;             
wire            clk_div_rst;             
wire            load_cmd;                
wire    [31:0]  m_haddr;                 
wire    [31:0]  m_haddr_fifo;            
wire    [31:0]  m_haddr_sub;             
wire    [2 :0]  m_hburst;                
wire    [2 :0]  m_hburst_fifo;           
wire    [2 :0]  m_hburst_sub;            
wire    [3 :0]  m_hprot;                 
wire    [3 :0]  m_hprot_fifo;            
wire    [3 :0]  m_hprot_sub;             
wire    [31:0]  m_hrdata;                
wire    [31:0]  m_hrdata_fifo;           
wire    [31:0]  m_hrdata_sub;            
wire            m_hready;                
wire            m_hready_fifo;           
wire            m_hready_sub;            
wire    [1 :0]  m_hresp;                 
wire    [1 :0]  m_hresp_fifo;            
wire    [1 :0]  m_hresp_sub;             
wire            m_hselx;                 
wire    [2 :0]  m_hsize;                 
wire    [2 :0]  m_hsize_fifo;            
wire    [2 :0]  m_hsize_sub;             
wire    [1 :0]  m_htrans;                
wire    [1 :0]  m_htrans_fifo;           
wire    [1 :0]  m_htrans_sub;            
wire    [31:0]  m_hwdata;                
wire    [31:0]  m_hwdata_fifo;           
wire    [31:0]  m_hwdata_sub;            
wire            m_hwrite;                
wire            m_hwrite_fifo;           
wire            m_hwrite_sub;            
wire            m_resp_vld;              
wire            m_resp_vld_sub;          
wire            main_hclk;               
wire            main_hresetn;            
wire            pmu_matrix_clkdiv_bypass; 
wire            rfifo_rd_aempty;         
wire    [34:0]  rfifo_rd_data;           
wire            rfifo_rd_empty;          
wire            rfifo_rd_en;             
wire            rfifo_rd_reset;          
wire            rfifo_wr_afull;          
wire    [34:0]  rfifo_wr_data;           
wire            rfifo_wr_en;             
wire            rfifo_wr_full;           
wire            rfifo_wr_reset;          
wire    [31:0]  s0_haddr;                
wire    [2 :0]  s0_hburst;               
wire    [3 :0]  s0_hprot;                
wire    [31:0]  s0_hrdata;               
wire            s0_hready;               
wire    [1 :0]  s0_hresp;                
wire            s0_hselx;                
wire    [2 :0]  s0_hsize;                
wire    [1 :0]  s0_htrans;               
wire    [31:0]  s0_hwdata;               
wire            s0_hwrite;               
wire    [31:0]  s1_haddr;                
wire    [2 :0]  s1_hburst;               
wire    [3 :0]  s1_hprot;                
wire    [31:0]  s1_hrdata;               
wire            s1_hready;               
wire    [1 :0]  s1_hresp;                
wire            s1_hselx;                
wire    [2 :0]  s1_hsize;                
wire    [1 :0]  s1_htrans;               
wire    [31:0]  s1_hwdata;               
wire            s1_hwrite;               
wire    [31:0]  s2_haddr;                
wire    [2 :0]  s2_hburst;               
wire    [3 :0]  s2_hprot;                
wire    [31:0]  s2_hrdata;               
wire            s2_hready;               
wire    [1 :0]  s2_hresp;                
wire            s2_hselx;                
wire    [2 :0]  s2_hsize;                
wire    [1 :0]  s2_htrans;               
wire    [31:0]  s2_hwdata;               
wire            s2_hwrite;               
wire    [31:0]  s3_haddr;                
wire    [2 :0]  s3_hburst;               
wire    [3 :0]  s3_hprot;                
wire    [31:0]  s3_hrdata;               
wire            s3_hready;               
wire    [1 :0]  s3_hresp;                
wire            s3_hselx;                
wire    [2 :0]  s3_hsize;                
wire    [1 :0]  s3_htrans;               
wire    [31:0]  s3_hwdata;               
wire            s3_hwrite;               
wire    [31:0]  s4_haddr;                
wire    [2 :0]  s4_hburst;               
wire    [3 :0]  s4_hprot;                
wire    [31:0]  s4_hrdata;               
wire            s4_hready;               
wire    [1 :0]  s4_hresp;                
wire            s4_hselx;                
wire    [2 :0]  s4_hsize;                
wire    [1 :0]  s4_htrans;               
wire    [31:0]  s4_hwdata;               
wire            s4_hwrite;               
wire    [31:0]  s5_haddr;                
wire    [2 :0]  s5_hburst;               
wire    [3 :0]  s5_hprot;                
wire    [31:0]  s5_hrdata;               
wire            s5_hready;               
wire    [1 :0]  s5_hresp;                
wire            s5_hselx;                
wire    [2 :0]  s5_hsize;                
wire    [1 :0]  s5_htrans;               
wire    [31:0]  s5_hwdata;               
wire            s5_hwrite;               
wire            sub_hclk;                
wire            sub_hresetn;             
wire            wfifo_rd_aempty;         
wire    [76:0]  wfifo_rd_data;           
wire            wfifo_rd_empty;          
wire            wfifo_rd_en;             
wire            wfifo_rd_reset;          
wire            wfifo_wr_afull;          
wire    [76:0]  wfifo_wr_data;           
wire            wfifo_wr_full;           
wire            wfifo_wr_reset;          
ahb_matrix_1_6_sub_dec  x_matrix_sub_dec (
  .hclk                     (sub_hclk                ),
  .hresetn                  (sub_hresetn             ),
  .load_cmd                 (load_cmd                ),
  .m_haddr                  (m_haddr_sub             ),
  .m_hburst                 (m_hburst_sub            ),
  .m_hprot                  (m_hprot_sub             ),
  .m_hrdata                 (m_hrdata_sub            ),
  .m_hready                 (m_hready_sub            ),
  .m_hresp                  (m_hresp_sub             ),
  .m_hsize                  (m_hsize_sub             ),
  .m_htrans                 (m_htrans_sub            ),
  .m_hwdata                 (m_hwdata_sub            ),
  .m_hwrite                 (m_hwrite_sub            ),
  .m_resp_vld               (m_resp_vld_sub          ),
  .pmu_matrix_clkdiv_bypass (pmu_matrix_clkdiv_bypass),
  .s0_haddr                 (s0_haddr                ),
  .s0_hburst                (s0_hburst               ),
  .s0_hprot                 (s0_hprot                ),
  .s0_hrdata                (s0_hrdata               ),
  .s0_hready                (s0_hready               ),
  .s0_hresp                 (s0_hresp                ),
  .s0_hselx                 (s0_hselx                ),
  .s0_hsize                 (s0_hsize                ),
  .s0_htrans                (s0_htrans               ),
  .s0_hwdata                (s0_hwdata               ),
  .s0_hwrite                (s0_hwrite               ),
  .s1_haddr                 (s1_haddr                ),
  .s1_hburst                (s1_hburst               ),
  .s1_hprot                 (s1_hprot                ),
  .s1_hrdata                (s1_hrdata               ),
  .s1_hready                (s1_hready               ),
  .s1_hresp                 (s1_hresp                ),
  .s1_hselx                 (s1_hselx                ),
  .s1_hsize                 (s1_hsize                ),
  .s1_htrans                (s1_htrans               ),
  .s1_hwdata                (s1_hwdata               ),
  .s1_hwrite                (s1_hwrite               ),
  .s2_haddr                 (s2_haddr                ),
  .s2_hburst                (s2_hburst               ),
  .s2_hprot                 (s2_hprot                ),
  .s2_hrdata                (s2_hrdata               ),
  .s2_hready                (s2_hready               ),
  .s2_hresp                 (s2_hresp                ),
  .s2_hselx                 (s2_hselx                ),
  .s2_hsize                 (s2_hsize                ),
  .s2_htrans                (s2_htrans               ),
  .s2_hwdata                (s2_hwdata               ),
  .s2_hwrite                (s2_hwrite               ),
  .s3_haddr                 (s3_haddr                ),
  .s3_hburst                (s3_hburst               ),
  .s3_hprot                 (s3_hprot                ),
  .s3_hrdata                (s3_hrdata               ),
  .s3_hready                (s3_hready               ),
  .s3_hresp                 (s3_hresp                ),
  .s3_hselx                 (s3_hselx                ),
  .s3_hsize                 (s3_hsize                ),
  .s3_htrans                (s3_htrans               ),
  .s3_hwdata                (s3_hwdata               ),
  .s3_hwrite                (s3_hwrite               ),
  .s4_haddr                 (s4_haddr                ),
  .s4_hburst                (s4_hburst               ),
  .s4_hprot                 (s4_hprot                ),
  .s4_hrdata                (s4_hrdata               ),
  .s4_hready                (s4_hready               ),
  .s4_hresp                 (s4_hresp                ),
  .s4_hselx                 (s4_hselx                ),
  .s4_hsize                 (s4_hsize                ),
  .s4_htrans                (s4_htrans               ),
  .s4_hwdata                (s4_hwdata               ),
  .s4_hwrite                (s4_hwrite               ),
  .s5_haddr                 (s5_haddr                ),
  .s5_hburst                (s5_hburst               ),
  .s5_hprot                 (s5_hprot                ),
  .s5_hrdata                (s5_hrdata               ),
  .s5_hready                (s5_hready               ),
  .s5_hresp                 (s5_hresp                ),
  .s5_hselx                 (s5_hselx                ),
  .s5_hsize                 (s5_hsize                ),
  .s5_htrans                (s5_htrans               ),
  .s5_hwdata                (s5_hwdata               ),
  .s5_hwrite                (s5_hwrite               ),
  .wfifo_rd_empty           (wfifo_rd_empty          )
);
afifo_77x2  x_sub_wr_afifo (
  .rd_aempty       (wfifo_rd_aempty),
  .rd_clk          (sub_hclk       ),
  .rd_data         (wfifo_rd_data  ),
  .rd_empty        (wfifo_rd_empty ),
  .rd_en           (wfifo_rd_en    ),
  .rd_reset_n      (wfifo_rd_reset ),
  .wr_afull        (wfifo_wr_afull ),
  .wr_clk          (main_hclk      ),
  .wr_data         (wfifo_wr_data  ),
  .wr_en           (wfifo_wr_en    ),
  .wr_full         (wfifo_wr_full  ),
  .wr_reset_n      (wfifo_wr_reset )
);
assign wfifo_wr_reset = main_hresetn & clk_div_rst;
assign wfifo_rd_reset = sub_hresetn & clk_div_rst;
always @ (posedge main_hclk or negedge main_hresetn)
    begin
       if(~main_hresetn)
         wfifo_wr_en <= 1'b0;
       else
         wfifo_wr_en <= ~wfifo_wr_afull & m_hselx & (~pmu_matrix_clkdiv_bypass);
    end
always @ (posedge main_hclk)
    begin
      m_haddr_d[31:0] <= m_haddr[31:0];
      m_htrans_d[1:0] <= m_htrans[1:0];
      m_hsize_d[2:0] <= m_hsize[2:0];
      m_hburst_d[2:0] <= m_hburst[2:0];
      m_hprot_d[3:0] <= m_hprot[3:0];
      m_hwrite_d <= m_hwrite;
    end
assign wfifo_wr_data[76:0] = {m_haddr_d[31:0],m_htrans_d[1:0],m_hsize_d[2:0],m_hburst_d[2:0],m_hprot_d[3:0],m_hwrite_d,m_hwdata[31:0]};
assign wfifo_rd_en = load_cmd;
assign {m_haddr_fifo[31:0],m_htrans_fifo[1:0],m_hsize_fifo[2:0],m_hburst_fifo[2:0],m_hprot_fifo[3:0],m_hwrite_fifo,m_hwdata_fifo[31:0]} = wfifo_rd_en ? wfifo_rd_data[76:0] : 77'd0;
afifo_35x2  x_sub_rd_afifo (
  .rd_aempty       (rfifo_rd_aempty),
  .rd_clk          (main_hclk      ),
  .rd_data         (rfifo_rd_data  ),
  .rd_empty        (rfifo_rd_empty ),
  .rd_en           (rfifo_rd_en    ),
  .rd_reset_n      (rfifo_rd_reset ),
  .wr_afull        (rfifo_wr_afull ),
  .wr_clk          (sub_hclk       ),
  .wr_data         (rfifo_wr_data  ),
  .wr_en           (rfifo_wr_en    ),
  .wr_full         (rfifo_wr_full  ),
  .wr_reset_n      (rfifo_wr_reset )
);
assign rfifo_wr_reset = sub_hresetn & clk_div_rst;
assign rfifo_rd_reset = main_hresetn & clk_div_rst;
assign rfifo_wr_en = (~rfifo_wr_afull) & m_resp_vld_sub & ~pmu_matrix_clkdiv_bypass;
assign rfifo_wr_data[34:0] = {m_hrdata_sub[31:0],m_hresp_sub[1:0],m_resp_vld_sub};
assign rfifo_rd_en = ~rfifo_rd_empty;
assign m_hrdata_fifo[31:0] = rfifo_rd_data[34:3];
assign m_hresp_fifo[1:0]= rfifo_rd_en ? rfifo_rd_data[2:1] : 2'b00;
assign m_resp_vld = rfifo_rd_en ? rfifo_rd_data[0] : 1'b0;
assign m_hready_fifo= (~wfifo_wr_full)&((~rd_hready)|m_resp_vld);
always @ (posedge main_hclk or negedge main_hresetn)
	begin
		if(~main_hresetn) begin
			rd_hready <= 1'b0;
		end
		else if(m_htrans[1]) begin
			rd_hready <= 1'b1;
		end
		else if(m_resp_vld) begin
			rd_hready <= 1'b0;
		end
	end
always @ (posedge main_hclk or negedge main_hresetn)
    begin
        if(~main_hresetn)
            clk_div <= 1'b0;
        else
            clk_div <= pmu_matrix_clkdiv_bypass;
    end
assign clk_div_rst = pmu_matrix_clkdiv_bypass | ~clk_div;
assign m_haddr_sub[31:0] = pmu_matrix_clkdiv_bypass ? m_haddr[31:0] : m_haddr_fifo[31:0];
assign m_htrans_sub[1:0] = pmu_matrix_clkdiv_bypass ? m_htrans[1:0] : m_htrans_fifo[1:0];
assign m_hburst_sub[2:0] = pmu_matrix_clkdiv_bypass ? m_hburst[2:0] : m_hburst_fifo[2:0];
assign m_hsize_sub[2:0]  = pmu_matrix_clkdiv_bypass ? m_hsize[2:0] : m_hsize_fifo[2:0];
assign m_hprot_sub[3:0]  = pmu_matrix_clkdiv_bypass ? m_hprot[3:0] : m_hprot_fifo[3:0];
assign m_hwrite_sub      = pmu_matrix_clkdiv_bypass ? m_hwrite : m_hwrite_fifo;
assign m_hwdata_sub[31:0]= pmu_matrix_clkdiv_bypass ? m_hwdata[31:0] : m_hwdata_fifo[31:0];
assign m_hrdata[31:0]    = pmu_matrix_clkdiv_bypass ? m_hrdata_sub[31:0] : m_hrdata_fifo[31:0];
assign m_hresp[1:0]      = pmu_matrix_clkdiv_bypass ? m_hresp_sub[1:0] : m_hresp_fifo[1:0];
assign m_hready          = pmu_matrix_clkdiv_bypass ? m_hready_sub : m_hready_fifo;
endmodule
module ahb_matrix_7_12_arb(
  hclk,
  hresetn,
  m0_latch_cmd,
  m0_nor_hready,
  m0_s0_cmd_cur,
  m0_s0_cmd_last,
  m0_s0_data,
  m0_s0_req,
  m0_s10_cmd_cur,
  m0_s10_cmd_last,
  m0_s10_data,
  m0_s10_req,
  m0_s11_cmd_cur,
  m0_s11_cmd_last,
  m0_s11_data,
  m0_s11_req,
  m0_s1_cmd_cur,
  m0_s1_cmd_last,
  m0_s1_data,
  m0_s1_req,
  m0_s2_cmd_cur,
  m0_s2_cmd_last,
  m0_s2_data,
  m0_s2_req,
  m0_s3_cmd_cur,
  m0_s3_cmd_last,
  m0_s3_data,
  m0_s3_req,
  m0_s4_cmd_cur,
  m0_s4_cmd_last,
  m0_s4_data,
  m0_s4_req,
  m0_s5_cmd_cur,
  m0_s5_cmd_last,
  m0_s5_data,
  m0_s5_req,
  m0_s6_cmd_cur,
  m0_s6_cmd_last,
  m0_s6_data,
  m0_s6_req,
  m0_s7_cmd_cur,
  m0_s7_cmd_last,
  m0_s7_data,
  m0_s7_req,
  m0_s8_cmd_cur,
  m0_s8_cmd_last,
  m0_s8_data,
  m0_s8_req,
  m0_s9_cmd_cur,
  m0_s9_cmd_last,
  m0_s9_data,
  m0_s9_req,
  m1_latch_cmd,
  m1_nor_hready,
  m1_s0_cmd_cur,
  m1_s0_cmd_last,
  m1_s0_data,
  m1_s0_req,
  m1_s10_cmd_cur,
  m1_s10_cmd_last,
  m1_s10_data,
  m1_s10_req,
  m1_s11_cmd_cur,
  m1_s11_cmd_last,
  m1_s11_data,
  m1_s11_req,
  m1_s1_cmd_cur,
  m1_s1_cmd_last,
  m1_s1_data,
  m1_s1_req,
  m1_s2_cmd_cur,
  m1_s2_cmd_last,
  m1_s2_data,
  m1_s2_req,
  m1_s3_cmd_cur,
  m1_s3_cmd_last,
  m1_s3_data,
  m1_s3_req,
  m1_s4_cmd_cur,
  m1_s4_cmd_last,
  m1_s4_data,
  m1_s4_req,
  m1_s5_cmd_cur,
  m1_s5_cmd_last,
  m1_s5_data,
  m1_s5_req,
  m1_s6_cmd_cur,
  m1_s6_cmd_last,
  m1_s6_data,
  m1_s6_req,
  m1_s7_cmd_cur,
  m1_s7_cmd_last,
  m1_s7_data,
  m1_s7_req,
  m1_s8_cmd_cur,
  m1_s8_cmd_last,
  m1_s8_data,
  m1_s8_req,
  m1_s9_cmd_cur,
  m1_s9_cmd_last,
  m1_s9_data,
  m1_s9_req,
  m2_latch_cmd,
  m2_nor_hready,
  m2_s0_cmd_cur,
  m2_s0_cmd_last,
  m2_s0_data,
  m2_s0_req,
  m2_s10_cmd_cur,
  m2_s10_cmd_last,
  m2_s10_data,
  m2_s10_req,
  m2_s11_cmd_cur,
  m2_s11_cmd_last,
  m2_s11_data,
  m2_s11_req,
  m2_s1_cmd_cur,
  m2_s1_cmd_last,
  m2_s1_data,
  m2_s1_req,
  m2_s2_cmd_cur,
  m2_s2_cmd_last,
  m2_s2_data,
  m2_s2_req,
  m2_s3_cmd_cur,
  m2_s3_cmd_last,
  m2_s3_data,
  m2_s3_req,
  m2_s4_cmd_cur,
  m2_s4_cmd_last,
  m2_s4_data,
  m2_s4_req,
  m2_s5_cmd_cur,
  m2_s5_cmd_last,
  m2_s5_data,
  m2_s5_req,
  m2_s6_cmd_cur,
  m2_s6_cmd_last,
  m2_s6_data,
  m2_s6_req,
  m2_s7_cmd_cur,
  m2_s7_cmd_last,
  m2_s7_data,
  m2_s7_req,
  m2_s8_cmd_cur,
  m2_s8_cmd_last,
  m2_s8_data,
  m2_s8_req,
  m2_s9_cmd_cur,
  m2_s9_cmd_last,
  m2_s9_data,
  m2_s9_req,
  m3_latch_cmd,
  m3_nor_hready,
  m3_s0_cmd_cur,
  m3_s0_cmd_last,
  m3_s0_data,
  m3_s0_req,
  m3_s10_cmd_cur,
  m3_s10_cmd_last,
  m3_s10_data,
  m3_s10_req,
  m3_s11_cmd_cur,
  m3_s11_cmd_last,
  m3_s11_data,
  m3_s11_req,
  m3_s1_cmd_cur,
  m3_s1_cmd_last,
  m3_s1_data,
  m3_s1_req,
  m3_s2_cmd_cur,
  m3_s2_cmd_last,
  m3_s2_data,
  m3_s2_req,
  m3_s3_cmd_cur,
  m3_s3_cmd_last,
  m3_s3_data,
  m3_s3_req,
  m3_s4_cmd_cur,
  m3_s4_cmd_last,
  m3_s4_data,
  m3_s4_req,
  m3_s5_cmd_cur,
  m3_s5_cmd_last,
  m3_s5_data,
  m3_s5_req,
  m3_s6_cmd_cur,
  m3_s6_cmd_last,
  m3_s6_data,
  m3_s6_req,
  m3_s7_cmd_cur,
  m3_s7_cmd_last,
  m3_s7_data,
  m3_s7_req,
  m3_s8_cmd_cur,
  m3_s8_cmd_last,
  m3_s8_data,
  m3_s8_req,
  m3_s9_cmd_cur,
  m3_s9_cmd_last,
  m3_s9_data,
  m3_s9_req,
  m4_latch_cmd,
  m4_nor_hready,
  m4_s0_cmd_cur,
  m4_s0_cmd_last,
  m4_s0_data,
  m4_s0_req,
  m4_s10_cmd_cur,
  m4_s10_cmd_last,
  m4_s10_data,
  m4_s10_req,
  m4_s11_cmd_cur,
  m4_s11_cmd_last,
  m4_s11_data,
  m4_s11_req,
  m4_s1_cmd_cur,
  m4_s1_cmd_last,
  m4_s1_data,
  m4_s1_req,
  m4_s2_cmd_cur,
  m4_s2_cmd_last,
  m4_s2_data,
  m4_s2_req,
  m4_s3_cmd_cur,
  m4_s3_cmd_last,
  m4_s3_data,
  m4_s3_req,
  m4_s4_cmd_cur,
  m4_s4_cmd_last,
  m4_s4_data,
  m4_s4_req,
  m4_s5_cmd_cur,
  m4_s5_cmd_last,
  m4_s5_data,
  m4_s5_req,
  m4_s6_cmd_cur,
  m4_s6_cmd_last,
  m4_s6_data,
  m4_s6_req,
  m4_s7_cmd_cur,
  m4_s7_cmd_last,
  m4_s7_data,
  m4_s7_req,
  m4_s8_cmd_cur,
  m4_s8_cmd_last,
  m4_s8_data,
  m4_s8_req,
  m4_s9_cmd_cur,
  m4_s9_cmd_last,
  m4_s9_data,
  m4_s9_req,
  m5_latch_cmd,
  m5_nor_hready,
  m5_s0_cmd_cur,
  m5_s0_cmd_last,
  m5_s0_data,
  m5_s0_req,
  m5_s10_cmd_cur,
  m5_s10_cmd_last,
  m5_s10_data,
  m5_s10_req,
  m5_s11_cmd_cur,
  m5_s11_cmd_last,
  m5_s11_data,
  m5_s11_req,
  m5_s1_cmd_cur,
  m5_s1_cmd_last,
  m5_s1_data,
  m5_s1_req,
  m5_s2_cmd_cur,
  m5_s2_cmd_last,
  m5_s2_data,
  m5_s2_req,
  m5_s3_cmd_cur,
  m5_s3_cmd_last,
  m5_s3_data,
  m5_s3_req,
  m5_s4_cmd_cur,
  m5_s4_cmd_last,
  m5_s4_data,
  m5_s4_req,
  m5_s5_cmd_cur,
  m5_s5_cmd_last,
  m5_s5_data,
  m5_s5_req,
  m5_s6_cmd_cur,
  m5_s6_cmd_last,
  m5_s6_data,
  m5_s6_req,
  m5_s7_cmd_cur,
  m5_s7_cmd_last,
  m5_s7_data,
  m5_s7_req,
  m5_s8_cmd_cur,
  m5_s8_cmd_last,
  m5_s8_data,
  m5_s8_req,
  m5_s9_cmd_cur,
  m5_s9_cmd_last,
  m5_s9_data,
  m5_s9_req,
  m6_latch_cmd,
  m6_nor_hready,
  m6_s0_cmd_cur,
  m6_s0_cmd_last,
  m6_s0_data,
  m6_s0_req,
  m6_s10_cmd_cur,
  m6_s10_cmd_last,
  m6_s10_data,
  m6_s10_req,
  m6_s11_cmd_cur,
  m6_s11_cmd_last,
  m6_s11_data,
  m6_s11_req,
  m6_s1_cmd_cur,
  m6_s1_cmd_last,
  m6_s1_data,
  m6_s1_req,
  m6_s2_cmd_cur,
  m6_s2_cmd_last,
  m6_s2_data,
  m6_s2_req,
  m6_s3_cmd_cur,
  m6_s3_cmd_last,
  m6_s3_data,
  m6_s3_req,
  m6_s4_cmd_cur,
  m6_s4_cmd_last,
  m6_s4_data,
  m6_s4_req,
  m6_s5_cmd_cur,
  m6_s5_cmd_last,
  m6_s5_data,
  m6_s5_req,
  m6_s6_cmd_cur,
  m6_s6_cmd_last,
  m6_s6_data,
  m6_s6_req,
  m6_s7_cmd_cur,
  m6_s7_cmd_last,
  m6_s7_data,
  m6_s7_req,
  m6_s8_cmd_cur,
  m6_s8_cmd_last,
  m6_s8_data,
  m6_s8_req,
  m6_s9_cmd_cur,
  m6_s9_cmd_last,
  m6_s9_data,
  m6_s9_req,
  s0_hready,
  s0_req,
  s10_hready,
  s10_req,
  s11_hready,
  s11_req,
  s1_hready,
  s1_req,
  s2_hready,
  s2_req,
  s3_hready,
  s3_req,
  s4_hready,
  s4_req,
  s5_hready,
  s5_req,
  s6_hready,
  s6_req,
  s7_hready,
  s7_req,
  s8_hready,
  s8_req,
  s9_hready,
  s9_req
);
input           hclk;               
input           hresetn;            
input           m0_s0_req;          
input           m0_s10_req;         
input           m0_s11_req;         
input           m0_s1_req;          
input           m0_s2_req;          
input           m0_s3_req;          
input           m0_s4_req;          
input           m0_s5_req;          
input           m0_s6_req;          
input           m0_s7_req;          
input           m0_s8_req;          
input           m0_s9_req;          
input           m1_s0_req;          
input           m1_s10_req;         
input           m1_s11_req;         
input           m1_s1_req;          
input           m1_s2_req;          
input           m1_s3_req;          
input           m1_s4_req;          
input           m1_s5_req;          
input           m1_s6_req;          
input           m1_s7_req;          
input           m1_s8_req;          
input           m1_s9_req;          
input           m2_s0_req;          
input           m2_s10_req;         
input           m2_s11_req;         
input           m2_s1_req;          
input           m2_s2_req;          
input           m2_s3_req;          
input           m2_s4_req;          
input           m2_s5_req;          
input           m2_s6_req;          
input           m2_s7_req;          
input           m2_s8_req;          
input           m2_s9_req;          
input           m3_s0_req;          
input           m3_s10_req;         
input           m3_s11_req;         
input           m3_s1_req;          
input           m3_s2_req;          
input           m3_s3_req;          
input           m3_s4_req;          
input           m3_s5_req;          
input           m3_s6_req;          
input           m3_s7_req;          
input           m3_s8_req;          
input           m3_s9_req;          
input           m4_s0_req;          
input           m4_s10_req;         
input           m4_s11_req;         
input           m4_s1_req;          
input           m4_s2_req;          
input           m4_s3_req;          
input           m4_s4_req;          
input           m4_s5_req;          
input           m4_s6_req;          
input           m4_s7_req;          
input           m4_s8_req;          
input           m4_s9_req;          
input           m5_s0_req;          
input           m5_s10_req;         
input           m5_s11_req;         
input           m5_s1_req;          
input           m5_s2_req;          
input           m5_s3_req;          
input           m5_s4_req;          
input           m5_s5_req;          
input           m5_s6_req;          
input           m5_s7_req;          
input           m5_s8_req;          
input           m5_s9_req;          
input           m6_s0_req;          
input           m6_s10_req;         
input           m6_s11_req;         
input           m6_s1_req;          
input           m6_s2_req;          
input           m6_s3_req;          
input           m6_s4_req;          
input           m6_s5_req;          
input           m6_s6_req;          
input           m6_s7_req;          
input           m6_s8_req;          
input           m6_s9_req;          
input           s0_hready;          
input   [6 :0]  s0_req;             
input           s10_hready;         
input   [6 :0]  s10_req;            
input           s11_hready;         
input   [6 :0]  s11_req;            
input           s1_hready;          
input   [6 :0]  s1_req;             
input           s2_hready;          
input   [6 :0]  s2_req;             
input           s3_hready;          
input   [6 :0]  s3_req;             
input           s4_hready;          
input   [6 :0]  s4_req;             
input           s5_hready;          
input   [6 :0]  s5_req;             
input           s6_hready;          
input   [6 :0]  s6_req;             
input           s7_hready;          
input   [6 :0]  s7_req;             
input           s8_hready;          
input   [6 :0]  s8_req;             
input           s9_hready;          
input   [6 :0]  s9_req;             
output          m0_latch_cmd;       
output          m0_nor_hready;      
output          m0_s0_cmd_cur;      
output          m0_s0_cmd_last;     
output          m0_s0_data;         
output          m0_s10_cmd_cur;     
output          m0_s10_cmd_last;    
output          m0_s10_data;        
output          m0_s11_cmd_cur;     
output          m0_s11_cmd_last;    
output          m0_s11_data;        
output          m0_s1_cmd_cur;      
output          m0_s1_cmd_last;     
output          m0_s1_data;         
output          m0_s2_cmd_cur;      
output          m0_s2_cmd_last;     
output          m0_s2_data;         
output          m0_s3_cmd_cur;      
output          m0_s3_cmd_last;     
output          m0_s3_data;         
output          m0_s4_cmd_cur;      
output          m0_s4_cmd_last;     
output          m0_s4_data;         
output          m0_s5_cmd_cur;      
output          m0_s5_cmd_last;     
output          m0_s5_data;         
output          m0_s6_cmd_cur;      
output          m0_s6_cmd_last;     
output          m0_s6_data;         
output          m0_s7_cmd_cur;      
output          m0_s7_cmd_last;     
output          m0_s7_data;         
output          m0_s8_cmd_cur;      
output          m0_s8_cmd_last;     
output          m0_s8_data;         
output          m0_s9_cmd_cur;      
output          m0_s9_cmd_last;     
output          m0_s9_data;         
output          m1_latch_cmd;       
output          m1_nor_hready;      
output          m1_s0_cmd_cur;      
output          m1_s0_cmd_last;     
output          m1_s0_data;         
output          m1_s10_cmd_cur;     
output          m1_s10_cmd_last;    
output          m1_s10_data;        
output          m1_s11_cmd_cur;     
output          m1_s11_cmd_last;    
output          m1_s11_data;        
output          m1_s1_cmd_cur;      
output          m1_s1_cmd_last;     
output          m1_s1_data;         
output          m1_s2_cmd_cur;      
output          m1_s2_cmd_last;     
output          m1_s2_data;         
output          m1_s3_cmd_cur;      
output          m1_s3_cmd_last;     
output          m1_s3_data;         
output          m1_s4_cmd_cur;      
output          m1_s4_cmd_last;     
output          m1_s4_data;         
output          m1_s5_cmd_cur;      
output          m1_s5_cmd_last;     
output          m1_s5_data;         
output          m1_s6_cmd_cur;      
output          m1_s6_cmd_last;     
output          m1_s6_data;         
output          m1_s7_cmd_cur;      
output          m1_s7_cmd_last;     
output          m1_s7_data;         
output          m1_s8_cmd_cur;      
output          m1_s8_cmd_last;     
output          m1_s8_data;         
output          m1_s9_cmd_cur;      
output          m1_s9_cmd_last;     
output          m1_s9_data;         
output          m2_latch_cmd;       
output          m2_nor_hready;      
output          m2_s0_cmd_cur;      
output          m2_s0_cmd_last;     
output          m2_s0_data;         
output          m2_s10_cmd_cur;     
output          m2_s10_cmd_last;    
output          m2_s10_data;        
output          m2_s11_cmd_cur;     
output          m2_s11_cmd_last;    
output          m2_s11_data;        
output          m2_s1_cmd_cur;      
output          m2_s1_cmd_last;     
output          m2_s1_data;         
output          m2_s2_cmd_cur;      
output          m2_s2_cmd_last;     
output          m2_s2_data;         
output          m2_s3_cmd_cur;      
output          m2_s3_cmd_last;     
output          m2_s3_data;         
output          m2_s4_cmd_cur;      
output          m2_s4_cmd_last;     
output          m2_s4_data;         
output          m2_s5_cmd_cur;      
output          m2_s5_cmd_last;     
output          m2_s5_data;         
output          m2_s6_cmd_cur;      
output          m2_s6_cmd_last;     
output          m2_s6_data;         
output          m2_s7_cmd_cur;      
output          m2_s7_cmd_last;     
output          m2_s7_data;         
output          m2_s8_cmd_cur;      
output          m2_s8_cmd_last;     
output          m2_s8_data;         
output          m2_s9_cmd_cur;      
output          m2_s9_cmd_last;     
output          m2_s9_data;         
output          m3_latch_cmd;       
output          m3_nor_hready;      
output          m3_s0_cmd_cur;      
output          m3_s0_cmd_last;     
output          m3_s0_data;         
output          m3_s10_cmd_cur;     
output          m3_s10_cmd_last;    
output          m3_s10_data;        
output          m3_s11_cmd_cur;     
output          m3_s11_cmd_last;    
output          m3_s11_data;        
output          m3_s1_cmd_cur;      
output          m3_s1_cmd_last;     
output          m3_s1_data;         
output          m3_s2_cmd_cur;      
output          m3_s2_cmd_last;     
output          m3_s2_data;         
output          m3_s3_cmd_cur;      
output          m3_s3_cmd_last;     
output          m3_s3_data;         
output          m3_s4_cmd_cur;      
output          m3_s4_cmd_last;     
output          m3_s4_data;         
output          m3_s5_cmd_cur;      
output          m3_s5_cmd_last;     
output          m3_s5_data;         
output          m3_s6_cmd_cur;      
output          m3_s6_cmd_last;     
output          m3_s6_data;         
output          m3_s7_cmd_cur;      
output          m3_s7_cmd_last;     
output          m3_s7_data;         
output          m3_s8_cmd_cur;      
output          m3_s8_cmd_last;     
output          m3_s8_data;         
output          m3_s9_cmd_cur;      
output          m3_s9_cmd_last;     
output          m3_s9_data;         
output          m4_latch_cmd;       
output          m4_nor_hready;      
output          m4_s0_cmd_cur;      
output          m4_s0_cmd_last;     
output          m4_s0_data;         
output          m4_s10_cmd_cur;     
output          m4_s10_cmd_last;    
output          m4_s10_data;        
output          m4_s11_cmd_cur;     
output          m4_s11_cmd_last;    
output          m4_s11_data;        
output          m4_s1_cmd_cur;      
output          m4_s1_cmd_last;     
output          m4_s1_data;         
output          m4_s2_cmd_cur;      
output          m4_s2_cmd_last;     
output          m4_s2_data;         
output          m4_s3_cmd_cur;      
output          m4_s3_cmd_last;     
output          m4_s3_data;         
output          m4_s4_cmd_cur;      
output          m4_s4_cmd_last;     
output          m4_s4_data;         
output          m4_s5_cmd_cur;      
output          m4_s5_cmd_last;     
output          m4_s5_data;         
output          m4_s6_cmd_cur;      
output          m4_s6_cmd_last;     
output          m4_s6_data;         
output          m4_s7_cmd_cur;      
output          m4_s7_cmd_last;     
output          m4_s7_data;         
output          m4_s8_cmd_cur;      
output          m4_s8_cmd_last;     
output          m4_s8_data;         
output          m4_s9_cmd_cur;      
output          m4_s9_cmd_last;     
output          m4_s9_data;         
output          m5_latch_cmd;       
output          m5_nor_hready;      
output          m5_s0_cmd_cur;      
output          m5_s0_cmd_last;     
output          m5_s0_data;         
output          m5_s10_cmd_cur;     
output          m5_s10_cmd_last;    
output          m5_s10_data;        
output          m5_s11_cmd_cur;     
output          m5_s11_cmd_last;    
output          m5_s11_data;        
output          m5_s1_cmd_cur;      
output          m5_s1_cmd_last;     
output          m5_s1_data;         
output          m5_s2_cmd_cur;      
output          m5_s2_cmd_last;     
output          m5_s2_data;         
output          m5_s3_cmd_cur;      
output          m5_s3_cmd_last;     
output          m5_s3_data;         
output          m5_s4_cmd_cur;      
output          m5_s4_cmd_last;     
output          m5_s4_data;         
output          m5_s5_cmd_cur;      
output          m5_s5_cmd_last;     
output          m5_s5_data;         
output          m5_s6_cmd_cur;      
output          m5_s6_cmd_last;     
output          m5_s6_data;         
output          m5_s7_cmd_cur;      
output          m5_s7_cmd_last;     
output          m5_s7_data;         
output          m5_s8_cmd_cur;      
output          m5_s8_cmd_last;     
output          m5_s8_data;         
output          m5_s9_cmd_cur;      
output          m5_s9_cmd_last;     
output          m5_s9_data;         
output          m6_latch_cmd;       
output          m6_nor_hready;      
output          m6_s0_cmd_cur;      
output          m6_s0_cmd_last;     
output          m6_s0_data;         
output          m6_s10_cmd_cur;     
output          m6_s10_cmd_last;    
output          m6_s10_data;        
output          m6_s11_cmd_cur;     
output          m6_s11_cmd_last;    
output          m6_s11_data;        
output          m6_s1_cmd_cur;      
output          m6_s1_cmd_last;     
output          m6_s1_data;         
output          m6_s2_cmd_cur;      
output          m6_s2_cmd_last;     
output          m6_s2_data;         
output          m6_s3_cmd_cur;      
output          m6_s3_cmd_last;     
output          m6_s3_data;         
output          m6_s4_cmd_cur;      
output          m6_s4_cmd_last;     
output          m6_s4_data;         
output          m6_s5_cmd_cur;      
output          m6_s5_cmd_last;     
output          m6_s5_data;         
output          m6_s6_cmd_cur;      
output          m6_s6_cmd_last;     
output          m6_s6_data;         
output          m6_s7_cmd_cur;      
output          m6_s7_cmd_last;     
output          m6_s7_data;         
output          m6_s8_cmd_cur;      
output          m6_s8_cmd_last;     
output          m6_s8_data;         
output          m6_s9_cmd_cur;      
output          m6_s9_cmd_last;     
output          m6_s9_data;         
reg     [48:0]  m0_cur_st;          
reg             m0_latch_cmd;       
reg             m0_nor_hready;      
reg     [48:0]  m0_nxt_st;          
reg             m0_s0_cmd_cur;      
reg             m0_s0_cmd_last;     
reg             m0_s0_data;         
reg             m0_s0_req_pend_tmp; 
reg             m0_s10_cmd_cur;     
reg             m0_s10_cmd_last;    
reg             m0_s10_data;        
reg             m0_s10_req_pend_tmp; 
reg             m0_s11_cmd_cur;     
reg             m0_s11_cmd_last;    
reg             m0_s11_data;        
reg             m0_s11_req_pend_tmp; 
reg             m0_s1_cmd_cur;      
reg             m0_s1_cmd_last;     
reg             m0_s1_data;         
reg             m0_s1_req_pend_tmp; 
reg             m0_s2_cmd_cur;      
reg             m0_s2_cmd_last;     
reg             m0_s2_data;         
reg             m0_s2_req_pend_tmp; 
reg             m0_s3_cmd_cur;      
reg             m0_s3_cmd_last;     
reg             m0_s3_data;         
reg             m0_s3_req_pend_tmp; 
reg             m0_s4_cmd_cur;      
reg             m0_s4_cmd_last;     
reg             m0_s4_data;         
reg             m0_s4_req_pend_tmp; 
reg             m0_s5_cmd_cur;      
reg             m0_s5_cmd_last;     
reg             m0_s5_data;         
reg             m0_s5_req_pend_tmp; 
reg             m0_s6_cmd_cur;      
reg             m0_s6_cmd_last;     
reg             m0_s6_data;         
reg             m0_s6_req_pend_tmp; 
reg             m0_s7_cmd_cur;      
reg             m0_s7_cmd_last;     
reg             m0_s7_data;         
reg             m0_s7_req_pend_tmp; 
reg             m0_s8_cmd_cur;      
reg             m0_s8_cmd_last;     
reg             m0_s8_data;         
reg             m0_s8_req_pend_tmp; 
reg             m0_s9_cmd_cur;      
reg             m0_s9_cmd_last;     
reg             m0_s9_data;         
reg             m0_s9_req_pend_tmp; 
reg     [48:0]  m1_cur_st;          
reg             m1_latch_cmd;       
reg             m1_nor_hready;      
reg     [48:0]  m1_nxt_st;          
reg             m1_s0_cmd_cur;      
reg             m1_s0_cmd_last;     
reg             m1_s0_data;         
reg             m1_s0_req_pend_tmp; 
reg             m1_s10_cmd_cur;     
reg             m1_s10_cmd_last;    
reg             m1_s10_data;        
reg             m1_s10_req_pend_tmp; 
reg             m1_s11_cmd_cur;     
reg             m1_s11_cmd_last;    
reg             m1_s11_data;        
reg             m1_s11_req_pend_tmp; 
reg             m1_s1_cmd_cur;      
reg             m1_s1_cmd_last;     
reg             m1_s1_data;         
reg             m1_s1_req_pend_tmp; 
reg             m1_s2_cmd_cur;      
reg             m1_s2_cmd_last;     
reg             m1_s2_data;         
reg             m1_s2_req_pend_tmp; 
reg             m1_s3_cmd_cur;      
reg             m1_s3_cmd_last;     
reg             m1_s3_data;         
reg             m1_s3_req_pend_tmp; 
reg             m1_s4_cmd_cur;      
reg             m1_s4_cmd_last;     
reg             m1_s4_data;         
reg             m1_s4_req_pend_tmp; 
reg             m1_s5_cmd_cur;      
reg             m1_s5_cmd_last;     
reg             m1_s5_data;         
reg             m1_s5_req_pend_tmp; 
reg             m1_s6_cmd_cur;      
reg             m1_s6_cmd_last;     
reg             m1_s6_data;         
reg             m1_s6_req_pend_tmp; 
reg             m1_s7_cmd_cur;      
reg             m1_s7_cmd_last;     
reg             m1_s7_data;         
reg             m1_s7_req_pend_tmp; 
reg             m1_s8_cmd_cur;      
reg             m1_s8_cmd_last;     
reg             m1_s8_data;         
reg             m1_s8_req_pend_tmp; 
reg             m1_s9_cmd_cur;      
reg             m1_s9_cmd_last;     
reg             m1_s9_data;         
reg             m1_s9_req_pend_tmp; 
reg     [48:0]  m2_cur_st;          
reg             m2_latch_cmd;       
reg             m2_nor_hready;      
reg     [48:0]  m2_nxt_st;          
reg             m2_s0_cmd_cur;      
reg             m2_s0_cmd_last;     
reg             m2_s0_data;         
reg             m2_s0_req_pend_tmp; 
reg             m2_s10_cmd_cur;     
reg             m2_s10_cmd_last;    
reg             m2_s10_data;        
reg             m2_s10_req_pend_tmp; 
reg             m2_s11_cmd_cur;     
reg             m2_s11_cmd_last;    
reg             m2_s11_data;        
reg             m2_s11_req_pend_tmp; 
reg             m2_s1_cmd_cur;      
reg             m2_s1_cmd_last;     
reg             m2_s1_data;         
reg             m2_s1_req_pend_tmp; 
reg             m2_s2_cmd_cur;      
reg             m2_s2_cmd_last;     
reg             m2_s2_data;         
reg             m2_s2_req_pend_tmp; 
reg             m2_s3_cmd_cur;      
reg             m2_s3_cmd_last;     
reg             m2_s3_data;         
reg             m2_s3_req_pend_tmp; 
reg             m2_s4_cmd_cur;      
reg             m2_s4_cmd_last;     
reg             m2_s4_data;         
reg             m2_s4_req_pend_tmp; 
reg             m2_s5_cmd_cur;      
reg             m2_s5_cmd_last;     
reg             m2_s5_data;         
reg             m2_s5_req_pend_tmp; 
reg             m2_s6_cmd_cur;      
reg             m2_s6_cmd_last;     
reg             m2_s6_data;         
reg             m2_s6_req_pend_tmp; 
reg             m2_s7_cmd_cur;      
reg             m2_s7_cmd_last;     
reg             m2_s7_data;         
reg             m2_s7_req_pend_tmp; 
reg             m2_s8_cmd_cur;      
reg             m2_s8_cmd_last;     
reg             m2_s8_data;         
reg             m2_s8_req_pend_tmp; 
reg             m2_s9_cmd_cur;      
reg             m2_s9_cmd_last;     
reg             m2_s9_data;         
reg             m2_s9_req_pend_tmp; 
reg     [48:0]  m3_cur_st;          
reg             m3_latch_cmd;       
reg             m3_nor_hready;      
reg     [48:0]  m3_nxt_st;          
reg             m3_s0_cmd_cur;      
reg             m3_s0_cmd_last;     
reg             m3_s0_data;         
reg             m3_s0_req_pend_tmp; 
reg             m3_s10_cmd_cur;     
reg             m3_s10_cmd_last;    
reg             m3_s10_data;        
reg             m3_s10_req_pend_tmp; 
reg             m3_s11_cmd_cur;     
reg             m3_s11_cmd_last;    
reg             m3_s11_data;        
reg             m3_s11_req_pend_tmp; 
reg             m3_s1_cmd_cur;      
reg             m3_s1_cmd_last;     
reg             m3_s1_data;         
reg             m3_s1_req_pend_tmp; 
reg             m3_s2_cmd_cur;      
reg             m3_s2_cmd_last;     
reg             m3_s2_data;         
reg             m3_s2_req_pend_tmp; 
reg             m3_s3_cmd_cur;      
reg             m3_s3_cmd_last;     
reg             m3_s3_data;         
reg             m3_s3_req_pend_tmp; 
reg             m3_s4_cmd_cur;      
reg             m3_s4_cmd_last;     
reg             m3_s4_data;         
reg             m3_s4_req_pend_tmp; 
reg             m3_s5_cmd_cur;      
reg             m3_s5_cmd_last;     
reg             m3_s5_data;         
reg             m3_s5_req_pend_tmp; 
reg             m3_s6_cmd_cur;      
reg             m3_s6_cmd_last;     
reg             m3_s6_data;         
reg             m3_s6_req_pend_tmp; 
reg             m3_s7_cmd_cur;      
reg             m3_s7_cmd_last;     
reg             m3_s7_data;         
reg             m3_s7_req_pend_tmp; 
reg             m3_s8_cmd_cur;      
reg             m3_s8_cmd_last;     
reg             m3_s8_data;         
reg             m3_s8_req_pend_tmp; 
reg             m3_s9_cmd_cur;      
reg             m3_s9_cmd_last;     
reg             m3_s9_data;         
reg             m3_s9_req_pend_tmp; 
reg     [48:0]  m4_cur_st;          
reg             m4_latch_cmd;       
reg             m4_nor_hready;      
reg     [48:0]  m4_nxt_st;          
reg             m4_s0_cmd_cur;      
reg             m4_s0_cmd_last;     
reg             m4_s0_data;         
reg             m4_s0_req_pend_tmp; 
reg             m4_s10_cmd_cur;     
reg             m4_s10_cmd_last;    
reg             m4_s10_data;        
reg             m4_s10_req_pend_tmp; 
reg             m4_s11_cmd_cur;     
reg             m4_s11_cmd_last;    
reg             m4_s11_data;        
reg             m4_s11_req_pend_tmp; 
reg             m4_s1_cmd_cur;      
reg             m4_s1_cmd_last;     
reg             m4_s1_data;         
reg             m4_s1_req_pend_tmp; 
reg             m4_s2_cmd_cur;      
reg             m4_s2_cmd_last;     
reg             m4_s2_data;         
reg             m4_s2_req_pend_tmp; 
reg             m4_s3_cmd_cur;      
reg             m4_s3_cmd_last;     
reg             m4_s3_data;         
reg             m4_s3_req_pend_tmp; 
reg             m4_s4_cmd_cur;      
reg             m4_s4_cmd_last;     
reg             m4_s4_data;         
reg             m4_s4_req_pend_tmp; 
reg             m4_s5_cmd_cur;      
reg             m4_s5_cmd_last;     
reg             m4_s5_data;         
reg             m4_s5_req_pend_tmp; 
reg             m4_s6_cmd_cur;      
reg             m4_s6_cmd_last;     
reg             m4_s6_data;         
reg             m4_s6_req_pend_tmp; 
reg             m4_s7_cmd_cur;      
reg             m4_s7_cmd_last;     
reg             m4_s7_data;         
reg             m4_s7_req_pend_tmp; 
reg             m4_s8_cmd_cur;      
reg             m4_s8_cmd_last;     
reg             m4_s8_data;         
reg             m4_s8_req_pend_tmp; 
reg             m4_s9_cmd_cur;      
reg             m4_s9_cmd_last;     
reg             m4_s9_data;         
reg             m4_s9_req_pend_tmp; 
reg     [48:0]  m5_cur_st;          
reg             m5_latch_cmd;       
reg             m5_nor_hready;      
reg     [48:0]  m5_nxt_st;          
reg             m5_s0_cmd_cur;      
reg             m5_s0_cmd_last;     
reg             m5_s0_data;         
reg             m5_s0_req_pend_tmp; 
reg             m5_s10_cmd_cur;     
reg             m5_s10_cmd_last;    
reg             m5_s10_data;        
reg             m5_s10_req_pend_tmp; 
reg             m5_s11_cmd_cur;     
reg             m5_s11_cmd_last;    
reg             m5_s11_data;        
reg             m5_s11_req_pend_tmp; 
reg             m5_s1_cmd_cur;      
reg             m5_s1_cmd_last;     
reg             m5_s1_data;         
reg             m5_s1_req_pend_tmp; 
reg             m5_s2_cmd_cur;      
reg             m5_s2_cmd_last;     
reg             m5_s2_data;         
reg             m5_s2_req_pend_tmp; 
reg             m5_s3_cmd_cur;      
reg             m5_s3_cmd_last;     
reg             m5_s3_data;         
reg             m5_s3_req_pend_tmp; 
reg             m5_s4_cmd_cur;      
reg             m5_s4_cmd_last;     
reg             m5_s4_data;         
reg             m5_s4_req_pend_tmp; 
reg             m5_s5_cmd_cur;      
reg             m5_s5_cmd_last;     
reg             m5_s5_data;         
reg             m5_s5_req_pend_tmp; 
reg             m5_s6_cmd_cur;      
reg             m5_s6_cmd_last;     
reg             m5_s6_data;         
reg             m5_s6_req_pend_tmp; 
reg             m5_s7_cmd_cur;      
reg             m5_s7_cmd_last;     
reg             m5_s7_data;         
reg             m5_s7_req_pend_tmp; 
reg             m5_s8_cmd_cur;      
reg             m5_s8_cmd_last;     
reg             m5_s8_data;         
reg             m5_s8_req_pend_tmp; 
reg             m5_s9_cmd_cur;      
reg             m5_s9_cmd_last;     
reg             m5_s9_data;         
reg             m5_s9_req_pend_tmp; 
reg     [48:0]  m6_cur_st;          
reg             m6_latch_cmd;       
reg             m6_nor_hready;      
reg     [48:0]  m6_nxt_st;          
reg             m6_s0_cmd_cur;      
reg             m6_s0_cmd_last;     
reg             m6_s0_data;         
reg             m6_s0_req_pend_tmp; 
reg             m6_s10_cmd_cur;     
reg             m6_s10_cmd_last;    
reg             m6_s10_data;        
reg             m6_s10_req_pend_tmp; 
reg             m6_s11_cmd_cur;     
reg             m6_s11_cmd_last;    
reg             m6_s11_data;        
reg             m6_s11_req_pend_tmp; 
reg             m6_s1_cmd_cur;      
reg             m6_s1_cmd_last;     
reg             m6_s1_data;         
reg             m6_s1_req_pend_tmp; 
reg             m6_s2_cmd_cur;      
reg             m6_s2_cmd_last;     
reg             m6_s2_data;         
reg             m6_s2_req_pend_tmp; 
reg             m6_s3_cmd_cur;      
reg             m6_s3_cmd_last;     
reg             m6_s3_data;         
reg             m6_s3_req_pend_tmp; 
reg             m6_s4_cmd_cur;      
reg             m6_s4_cmd_last;     
reg             m6_s4_data;         
reg             m6_s4_req_pend_tmp; 
reg             m6_s5_cmd_cur;      
reg             m6_s5_cmd_last;     
reg             m6_s5_data;         
reg             m6_s5_req_pend_tmp; 
reg             m6_s6_cmd_cur;      
reg             m6_s6_cmd_last;     
reg             m6_s6_data;         
reg             m6_s6_req_pend_tmp; 
reg             m6_s7_cmd_cur;      
reg             m6_s7_cmd_last;     
reg             m6_s7_data;         
reg             m6_s7_req_pend_tmp; 
reg             m6_s8_cmd_cur;      
reg             m6_s8_cmd_last;     
reg             m6_s8_data;         
reg             m6_s8_req_pend_tmp; 
reg             m6_s9_cmd_cur;      
reg             m6_s9_cmd_last;     
reg             m6_s9_data;         
reg             m6_s9_req_pend_tmp; 
reg     [6 :0]  s0_gnt;             
reg     [6 :0]  s10_gnt;            
reg     [6 :0]  s11_gnt;            
reg     [6 :0]  s1_gnt;             
reg     [6 :0]  s2_gnt;             
reg     [6 :0]  s3_gnt;             
reg     [6 :0]  s4_gnt;             
reg     [6 :0]  s5_gnt;             
reg     [6 :0]  s6_gnt;             
reg     [6 :0]  s7_gnt;             
reg     [6 :0]  s8_gnt;             
reg     [6 :0]  s9_gnt;             
wire            hclk;               
wire            hresetn;            
wire            m0_s0_hld;          
wire            m0_s0_req;          
wire            m0_s0_req_pend;     
wire            m0_s0_sel;          
wire            m0_s0_wt_sel;       
wire            m0_s10_hld;         
wire            m0_s10_req;         
wire            m0_s10_req_pend;    
wire            m0_s10_sel;         
wire            m0_s10_wt_sel;      
wire            m0_s11_hld;         
wire            m0_s11_req;         
wire            m0_s11_req_pend;    
wire            m0_s11_sel;         
wire            m0_s11_wt_sel;      
wire            m0_s1_hld;          
wire            m0_s1_req;          
wire            m0_s1_req_pend;     
wire            m0_s1_sel;          
wire            m0_s1_wt_sel;       
wire            m0_s2_hld;          
wire            m0_s2_req;          
wire            m0_s2_req_pend;     
wire            m0_s2_sel;          
wire            m0_s2_wt_sel;       
wire            m0_s3_hld;          
wire            m0_s3_req;          
wire            m0_s3_req_pend;     
wire            m0_s3_sel;          
wire            m0_s3_wt_sel;       
wire            m0_s4_hld;          
wire            m0_s4_req;          
wire            m0_s4_req_pend;     
wire            m0_s4_sel;          
wire            m0_s4_wt_sel;       
wire            m0_s5_hld;          
wire            m0_s5_req;          
wire            m0_s5_req_pend;     
wire            m0_s5_sel;          
wire            m0_s5_wt_sel;       
wire            m0_s6_hld;          
wire            m0_s6_req;          
wire            m0_s6_req_pend;     
wire            m0_s6_sel;          
wire            m0_s6_wt_sel;       
wire            m0_s7_hld;          
wire            m0_s7_req;          
wire            m0_s7_req_pend;     
wire            m0_s7_sel;          
wire            m0_s7_wt_sel;       
wire            m0_s8_hld;          
wire            m0_s8_req;          
wire            m0_s8_req_pend;     
wire            m0_s8_sel;          
wire            m0_s8_wt_sel;       
wire            m0_s9_hld;          
wire            m0_s9_req;          
wire            m0_s9_req_pend;     
wire            m0_s9_sel;          
wire            m0_s9_wt_sel;       
wire            m1_s0_hld;          
wire            m1_s0_req;          
wire            m1_s0_req_pend;     
wire            m1_s0_sel;          
wire            m1_s0_wt_sel;       
wire            m1_s10_hld;         
wire            m1_s10_req;         
wire            m1_s10_req_pend;    
wire            m1_s10_sel;         
wire            m1_s10_wt_sel;      
wire            m1_s11_hld;         
wire            m1_s11_req;         
wire            m1_s11_req_pend;    
wire            m1_s11_sel;         
wire            m1_s11_wt_sel;      
wire            m1_s1_hld;          
wire            m1_s1_req;          
wire            m1_s1_req_pend;     
wire            m1_s1_sel;          
wire            m1_s1_wt_sel;       
wire            m1_s2_hld;          
wire            m1_s2_req;          
wire            m1_s2_req_pend;     
wire            m1_s2_sel;          
wire            m1_s2_wt_sel;       
wire            m1_s3_hld;          
wire            m1_s3_req;          
wire            m1_s3_req_pend;     
wire            m1_s3_sel;          
wire            m1_s3_wt_sel;       
wire            m1_s4_hld;          
wire            m1_s4_req;          
wire            m1_s4_req_pend;     
wire            m1_s4_sel;          
wire            m1_s4_wt_sel;       
wire            m1_s5_hld;          
wire            m1_s5_req;          
wire            m1_s5_req_pend;     
wire            m1_s5_sel;          
wire            m1_s5_wt_sel;       
wire            m1_s6_hld;          
wire            m1_s6_req;          
wire            m1_s6_req_pend;     
wire            m1_s6_sel;          
wire            m1_s6_wt_sel;       
wire            m1_s7_hld;          
wire            m1_s7_req;          
wire            m1_s7_req_pend;     
wire            m1_s7_sel;          
wire            m1_s7_wt_sel;       
wire            m1_s8_hld;          
wire            m1_s8_req;          
wire            m1_s8_req_pend;     
wire            m1_s8_sel;          
wire            m1_s8_wt_sel;       
wire            m1_s9_hld;          
wire            m1_s9_req;          
wire            m1_s9_req_pend;     
wire            m1_s9_sel;          
wire            m1_s9_wt_sel;       
wire            m2_s0_hld;          
wire            m2_s0_req;          
wire            m2_s0_req_pend;     
wire            m2_s0_sel;          
wire            m2_s0_wt_sel;       
wire            m2_s10_hld;         
wire            m2_s10_req;         
wire            m2_s10_req_pend;    
wire            m2_s10_sel;         
wire            m2_s10_wt_sel;      
wire            m2_s11_hld;         
wire            m2_s11_req;         
wire            m2_s11_req_pend;    
wire            m2_s11_sel;         
wire            m2_s11_wt_sel;      
wire            m2_s1_hld;          
wire            m2_s1_req;          
wire            m2_s1_req_pend;     
wire            m2_s1_sel;          
wire            m2_s1_wt_sel;       
wire            m2_s2_hld;          
wire            m2_s2_req;          
wire            m2_s2_req_pend;     
wire            m2_s2_sel;          
wire            m2_s2_wt_sel;       
wire            m2_s3_hld;          
wire            m2_s3_req;          
wire            m2_s3_req_pend;     
wire            m2_s3_sel;          
wire            m2_s3_wt_sel;       
wire            m2_s4_hld;          
wire            m2_s4_req;          
wire            m2_s4_req_pend;     
wire            m2_s4_sel;          
wire            m2_s4_wt_sel;       
wire            m2_s5_hld;          
wire            m2_s5_req;          
wire            m2_s5_req_pend;     
wire            m2_s5_sel;          
wire            m2_s5_wt_sel;       
wire            m2_s6_hld;          
wire            m2_s6_req;          
wire            m2_s6_req_pend;     
wire            m2_s6_sel;          
wire            m2_s6_wt_sel;       
wire            m2_s7_hld;          
wire            m2_s7_req;          
wire            m2_s7_req_pend;     
wire            m2_s7_sel;          
wire            m2_s7_wt_sel;       
wire            m2_s8_hld;          
wire            m2_s8_req;          
wire            m2_s8_req_pend;     
wire            m2_s8_sel;          
wire            m2_s8_wt_sel;       
wire            m2_s9_hld;          
wire            m2_s9_req;          
wire            m2_s9_req_pend;     
wire            m2_s9_sel;          
wire            m2_s9_wt_sel;       
wire            m3_s0_hld;          
wire            m3_s0_req;          
wire            m3_s0_req_pend;     
wire            m3_s0_sel;          
wire            m3_s0_wt_sel;       
wire            m3_s10_hld;         
wire            m3_s10_req;         
wire            m3_s10_req_pend;    
wire            m3_s10_sel;         
wire            m3_s10_wt_sel;      
wire            m3_s11_hld;         
wire            m3_s11_req;         
wire            m3_s11_req_pend;    
wire            m3_s11_sel;         
wire            m3_s11_wt_sel;      
wire            m3_s1_hld;          
wire            m3_s1_req;          
wire            m3_s1_req_pend;     
wire            m3_s1_sel;          
wire            m3_s1_wt_sel;       
wire            m3_s2_hld;          
wire            m3_s2_req;          
wire            m3_s2_req_pend;     
wire            m3_s2_sel;          
wire            m3_s2_wt_sel;       
wire            m3_s3_hld;          
wire            m3_s3_req;          
wire            m3_s3_req_pend;     
wire            m3_s3_sel;          
wire            m3_s3_wt_sel;       
wire            m3_s4_hld;          
wire            m3_s4_req;          
wire            m3_s4_req_pend;     
wire            m3_s4_sel;          
wire            m3_s4_wt_sel;       
wire            m3_s5_hld;          
wire            m3_s5_req;          
wire            m3_s5_req_pend;     
wire            m3_s5_sel;          
wire            m3_s5_wt_sel;       
wire            m3_s6_hld;          
wire            m3_s6_req;          
wire            m3_s6_req_pend;     
wire            m3_s6_sel;          
wire            m3_s6_wt_sel;       
wire            m3_s7_hld;          
wire            m3_s7_req;          
wire            m3_s7_req_pend;     
wire            m3_s7_sel;          
wire            m3_s7_wt_sel;       
wire            m3_s8_hld;          
wire            m3_s8_req;          
wire            m3_s8_req_pend;     
wire            m3_s8_sel;          
wire            m3_s8_wt_sel;       
wire            m3_s9_hld;          
wire            m3_s9_req;          
wire            m3_s9_req_pend;     
wire            m3_s9_sel;          
wire            m3_s9_wt_sel;       
wire            m4_s0_hld;          
wire            m4_s0_req;          
wire            m4_s0_req_pend;     
wire            m4_s0_sel;          
wire            m4_s0_wt_sel;       
wire            m4_s10_hld;         
wire            m4_s10_req;         
wire            m4_s10_req_pend;    
wire            m4_s10_sel;         
wire            m4_s10_wt_sel;      
wire            m4_s11_hld;         
wire            m4_s11_req;         
wire            m4_s11_req_pend;    
wire            m4_s11_sel;         
wire            m4_s11_wt_sel;      
wire            m4_s1_hld;          
wire            m4_s1_req;          
wire            m4_s1_req_pend;     
wire            m4_s1_sel;          
wire            m4_s1_wt_sel;       
wire            m4_s2_hld;          
wire            m4_s2_req;          
wire            m4_s2_req_pend;     
wire            m4_s2_sel;          
wire            m4_s2_wt_sel;       
wire            m4_s3_hld;          
wire            m4_s3_req;          
wire            m4_s3_req_pend;     
wire            m4_s3_sel;          
wire            m4_s3_wt_sel;       
wire            m4_s4_hld;          
wire            m4_s4_req;          
wire            m4_s4_req_pend;     
wire            m4_s4_sel;          
wire            m4_s4_wt_sel;       
wire            m4_s5_hld;          
wire            m4_s5_req;          
wire            m4_s5_req_pend;     
wire            m4_s5_sel;          
wire            m4_s5_wt_sel;       
wire            m4_s6_hld;          
wire            m4_s6_req;          
wire            m4_s6_req_pend;     
wire            m4_s6_sel;          
wire            m4_s6_wt_sel;       
wire            m4_s7_hld;          
wire            m4_s7_req;          
wire            m4_s7_req_pend;     
wire            m4_s7_sel;          
wire            m4_s7_wt_sel;       
wire            m4_s8_hld;          
wire            m4_s8_req;          
wire            m4_s8_req_pend;     
wire            m4_s8_sel;          
wire            m4_s8_wt_sel;       
wire            m4_s9_hld;          
wire            m4_s9_req;          
wire            m4_s9_req_pend;     
wire            m4_s9_sel;          
wire            m4_s9_wt_sel;       
wire            m5_s0_hld;          
wire            m5_s0_req;          
wire            m5_s0_req_pend;     
wire            m5_s0_sel;          
wire            m5_s0_wt_sel;       
wire            m5_s10_hld;         
wire            m5_s10_req;         
wire            m5_s10_req_pend;    
wire            m5_s10_sel;         
wire            m5_s10_wt_sel;      
wire            m5_s11_hld;         
wire            m5_s11_req;         
wire            m5_s11_req_pend;    
wire            m5_s11_sel;         
wire            m5_s11_wt_sel;      
wire            m5_s1_hld;          
wire            m5_s1_req;          
wire            m5_s1_req_pend;     
wire            m5_s1_sel;          
wire            m5_s1_wt_sel;       
wire            m5_s2_hld;          
wire            m5_s2_req;          
wire            m5_s2_req_pend;     
wire            m5_s2_sel;          
wire            m5_s2_wt_sel;       
wire            m5_s3_hld;          
wire            m5_s3_req;          
wire            m5_s3_req_pend;     
wire            m5_s3_sel;          
wire            m5_s3_wt_sel;       
wire            m5_s4_hld;          
wire            m5_s4_req;          
wire            m5_s4_req_pend;     
wire            m5_s4_sel;          
wire            m5_s4_wt_sel;       
wire            m5_s5_hld;          
wire            m5_s5_req;          
wire            m5_s5_req_pend;     
wire            m5_s5_sel;          
wire            m5_s5_wt_sel;       
wire            m5_s6_hld;          
wire            m5_s6_req;          
wire            m5_s6_req_pend;     
wire            m5_s6_sel;          
wire            m5_s6_wt_sel;       
wire            m5_s7_hld;          
wire            m5_s7_req;          
wire            m5_s7_req_pend;     
wire            m5_s7_sel;          
wire            m5_s7_wt_sel;       
wire            m5_s8_hld;          
wire            m5_s8_req;          
wire            m5_s8_req_pend;     
wire            m5_s8_sel;          
wire            m5_s8_wt_sel;       
wire            m5_s9_hld;          
wire            m5_s9_req;          
wire            m5_s9_req_pend;     
wire            m5_s9_sel;          
wire            m5_s9_wt_sel;       
wire            m6_s0_hld;          
wire            m6_s0_req;          
wire            m6_s0_req_pend;     
wire            m6_s0_sel;          
wire            m6_s0_wt_sel;       
wire            m6_s10_hld;         
wire            m6_s10_req;         
wire            m6_s10_req_pend;    
wire            m6_s10_sel;         
wire            m6_s10_wt_sel;      
wire            m6_s11_hld;         
wire            m6_s11_req;         
wire            m6_s11_req_pend;    
wire            m6_s11_sel;         
wire            m6_s11_wt_sel;      
wire            m6_s1_hld;          
wire            m6_s1_req;          
wire            m6_s1_req_pend;     
wire            m6_s1_sel;          
wire            m6_s1_wt_sel;       
wire            m6_s2_hld;          
wire            m6_s2_req;          
wire            m6_s2_req_pend;     
wire            m6_s2_sel;          
wire            m6_s2_wt_sel;       
wire            m6_s3_hld;          
wire            m6_s3_req;          
wire            m6_s3_req_pend;     
wire            m6_s3_sel;          
wire            m6_s3_wt_sel;       
wire            m6_s4_hld;          
wire            m6_s4_req;          
wire            m6_s4_req_pend;     
wire            m6_s4_sel;          
wire            m6_s4_wt_sel;       
wire            m6_s5_hld;          
wire            m6_s5_req;          
wire            m6_s5_req_pend;     
wire            m6_s5_sel;          
wire            m6_s5_wt_sel;       
wire            m6_s6_hld;          
wire            m6_s6_req;          
wire            m6_s6_req_pend;     
wire            m6_s6_sel;          
wire            m6_s6_wt_sel;       
wire            m6_s7_hld;          
wire            m6_s7_req;          
wire            m6_s7_req_pend;     
wire            m6_s7_sel;          
wire            m6_s7_wt_sel;       
wire            m6_s8_hld;          
wire            m6_s8_req;          
wire            m6_s8_req_pend;     
wire            m6_s8_sel;          
wire            m6_s8_wt_sel;       
wire            m6_s9_hld;          
wire            m6_s9_req;          
wire            m6_s9_req_pend;     
wire            m6_s9_sel;          
wire            m6_s9_wt_sel;       
wire            s0_hready;          
wire    [6 :0]  s0_req;             
wire    [6 :0]  s0_req_all;         
wire    [6 :0]  s0_req_pend;        
wire            s10_hready;         
wire    [6 :0]  s10_req;            
wire    [6 :0]  s10_req_all;        
wire    [6 :0]  s10_req_pend;       
wire            s11_hready;         
wire    [6 :0]  s11_req;            
wire    [6 :0]  s11_req_all;        
wire    [6 :0]  s11_req_pend;       
wire            s1_hready;          
wire    [6 :0]  s1_req;             
wire    [6 :0]  s1_req_all;         
wire    [6 :0]  s1_req_pend;        
wire            s2_hready;          
wire    [6 :0]  s2_req;             
wire    [6 :0]  s2_req_all;         
wire    [6 :0]  s2_req_pend;        
wire            s3_hready;          
wire    [6 :0]  s3_req;             
wire    [6 :0]  s3_req_all;         
wire    [6 :0]  s3_req_pend;        
wire            s4_hready;          
wire    [6 :0]  s4_req;             
wire    [6 :0]  s4_req_all;         
wire    [6 :0]  s4_req_pend;        
wire            s5_hready;          
wire    [6 :0]  s5_req;             
wire    [6 :0]  s5_req_all;         
wire    [6 :0]  s5_req_pend;        
wire            s6_hready;          
wire    [6 :0]  s6_req;             
wire    [6 :0]  s6_req_all;         
wire    [6 :0]  s6_req_pend;        
wire            s7_hready;          
wire    [6 :0]  s7_req;             
wire    [6 :0]  s7_req_all;         
wire    [6 :0]  s7_req_pend;        
wire            s8_hready;          
wire    [6 :0]  s8_req;             
wire    [6 :0]  s8_req_all;         
wire    [6 :0]  s8_req_pend;        
wire            s9_hready;          
wire    [6 :0]  s9_req;             
wire    [6 :0]  s9_req_all;         
wire    [6 :0]  s9_req_pend;        
parameter S_IDLE    = 49'b0000000000000000000000000000000000000000000000001;
parameter S_S0_GNT  = 49'b0000000000000000000000000000000000000000000000010;
parameter S_S0_WAIT = 49'b0000000000000000000000000000000000000000000000100;
parameter S_S0_CMD  = 49'b0000000000000000000000000000000000000000000001000;
parameter S_S0_DATA = 49'b0000000000000000000000000000000000000000000010000;
parameter S_S1_GNT  = 49'b0000000000000000000000000000000000000000000100000;
parameter S_S1_WAIT = 49'b0000000000000000000000000000000000000000001000000;
parameter S_S1_CMD  = 49'b0000000000000000000000000000000000000000010000000;
parameter S_S1_DATA = 49'b0000000000000000000000000000000000000000100000000;
parameter S_S2_GNT  = 49'b0000000000000000000000000000000000000001000000000;
parameter S_S2_WAIT = 49'b0000000000000000000000000000000000000010000000000;
parameter S_S2_CMD  = 49'b0000000000000000000000000000000000000100000000000;
parameter S_S2_DATA = 49'b0000000000000000000000000000000000001000000000000;
parameter S_S3_GNT  = 49'b0000000000000000000000000000000000010000000000000;
parameter S_S3_WAIT = 49'b0000000000000000000000000000000000100000000000000;
parameter S_S3_CMD  = 49'b0000000000000000000000000000000001000000000000000;
parameter S_S3_DATA = 49'b0000000000000000000000000000000010000000000000000;
parameter S_S4_GNT  = 49'b0000000000000000000000000000000100000000000000000;
parameter S_S4_WAIT = 49'b0000000000000000000000000000001000000000000000000;
parameter S_S4_CMD  = 49'b0000000000000000000000000000010000000000000000000;
parameter S_S4_DATA = 49'b0000000000000000000000000000100000000000000000000;
parameter S_S5_GNT  = 49'b0000000000000000000000000001000000000000000000000;
parameter S_S5_WAIT = 49'b0000000000000000000000000010000000000000000000000;
parameter S_S5_CMD  = 49'b0000000000000000000000000100000000000000000000000;
parameter S_S5_DATA = 49'b0000000000000000000000001000000000000000000000000;
parameter S_S6_GNT  = 49'b0000000000000000000000010000000000000000000000000;
parameter S_S6_WAIT = 49'b0000000000000000000000100000000000000000000000000;
parameter S_S6_CMD  = 49'b0000000000000000000001000000000000000000000000000;
parameter S_S6_DATA = 49'b0000000000000000000010000000000000000000000000000;
parameter S_S7_GNT  = 49'b0000000000000000000100000000000000000000000000000;
parameter S_S7_WAIT = 49'b0000000000000000001000000000000000000000000000000;
parameter S_S7_CMD  = 49'b0000000000000000010000000000000000000000000000000;
parameter S_S7_DATA = 49'b0000000000000000100000000000000000000000000000000;
parameter S_S8_GNT  = 49'b0000000000000001000000000000000000000000000000000;
parameter S_S8_WAIT = 49'b0000000000000010000000000000000000000000000000000;
parameter S_S8_CMD  = 49'b0000000000000100000000000000000000000000000000000;
parameter S_S8_DATA = 49'b0000000000001000000000000000000000000000000000000;
parameter S_S9_GNT  = 49'b0000000000010000000000000000000000000000000000000;
parameter S_S9_WAIT = 49'b0000000000100000000000000000000000000000000000000;
parameter S_S9_CMD  = 49'b0000000001000000000000000000000000000000000000000;
parameter S_S9_DATA = 49'b0000000010000000000000000000000000000000000000000;
parameter S_S10_GNT  = 49'b0000000100000000000000000000000000000000000000000;
parameter S_S10_WAIT = 49'b0000001000000000000000000000000000000000000000000;
parameter S_S10_CMD  = 49'b0000010000000000000000000000000000000000000000000;
parameter S_S10_DATA = 49'b0000100000000000000000000000000000000000000000000;
parameter S_S11_GNT  = 49'b0001000000000000000000000000000000000000000000000;
parameter S_S11_WAIT = 49'b0010000000000000000000000000000000000000000000000;
parameter S_S11_CMD  = 49'b0100000000000000000000000000000000000000000000000;
parameter S_S11_DATA = 49'b1000000000000000000000000000000000000000000000000;
assign s0_req_all[7-1:0] = s0_req[7-1:0] | s0_req_pend[7-1:0];
always @( s0_req_all[6:0])
begin
casez(s0_req_all[7-1:0])
   7'b1??????: s0_gnt[7-1:0] = 7'b1000000;
   7'b01?????: s0_gnt[7-1:0] = 7'b0100000;
   7'b001????: s0_gnt[7-1:0] = 7'b0010000;
   7'b0001???: s0_gnt[7-1:0] = 7'b0001000;
   7'b00001??: s0_gnt[7-1:0] = 7'b0000100;
   7'b000001?: s0_gnt[7-1:0] = 7'b0000010;
   7'b0000001: s0_gnt[7-1:0] = 7'b0000001;
   default: s0_gnt[7-1:0] = 7'b0000000;
endcase
end
assign s1_req_all[7-1:0] = s1_req[7-1:0] | s1_req_pend[7-1:0];
always @( s1_req_all[6:0])
begin
casez(s1_req_all[7-1:0])
   7'b1??????: s1_gnt[7-1:0] = 7'b1000000;
   7'b01?????: s1_gnt[7-1:0] = 7'b0100000;
   7'b001????: s1_gnt[7-1:0] = 7'b0010000;
   7'b0001???: s1_gnt[7-1:0] = 7'b0001000;
   7'b00001??: s1_gnt[7-1:0] = 7'b0000100;
   7'b000001?: s1_gnt[7-1:0] = 7'b0000010;
   7'b0000001: s1_gnt[7-1:0] = 7'b0000001;
   default: s1_gnt[7-1:0] = 7'b0000000;
endcase
end
assign s2_req_all[7-1:0] = s2_req[7-1:0] | s2_req_pend[7-1:0];
always @( s2_req_all[6:0])
begin
casez(s2_req_all[7-1:0])
   7'b1??????: s2_gnt[7-1:0] = 7'b1000000;
   7'b01?????: s2_gnt[7-1:0] = 7'b0100000;
   7'b001????: s2_gnt[7-1:0] = 7'b0010000;
   7'b0001???: s2_gnt[7-1:0] = 7'b0001000;
   7'b00001??: s2_gnt[7-1:0] = 7'b0000100;
   7'b000001?: s2_gnt[7-1:0] = 7'b0000010;
   7'b0000001: s2_gnt[7-1:0] = 7'b0000001;
   default: s2_gnt[7-1:0] = 7'b0000000;
endcase
end
assign s3_req_all[7-1:0] = s3_req[7-1:0] | s3_req_pend[7-1:0];
always @( s3_req_all[6:0])
begin
casez(s3_req_all[7-1:0])
   7'b1??????: s3_gnt[7-1:0] = 7'b1000000;
   7'b01?????: s3_gnt[7-1:0] = 7'b0100000;
   7'b001????: s3_gnt[7-1:0] = 7'b0010000;
   7'b0001???: s3_gnt[7-1:0] = 7'b0001000;
   7'b00001??: s3_gnt[7-1:0] = 7'b0000100;
   7'b000001?: s3_gnt[7-1:0] = 7'b0000010;
   7'b0000001: s3_gnt[7-1:0] = 7'b0000001;
   default: s3_gnt[7-1:0] = 7'b0000000;
endcase
end
assign s4_req_all[7-1:0] = s4_req[7-1:0] | s4_req_pend[7-1:0];
always @( s4_req_all[6:0])
begin
casez(s4_req_all[7-1:0])
   7'b1??????: s4_gnt[7-1:0] = 7'b1000000;
   7'b01?????: s4_gnt[7-1:0] = 7'b0100000;
   7'b001????: s4_gnt[7-1:0] = 7'b0010000;
   7'b0001???: s4_gnt[7-1:0] = 7'b0001000;
   7'b00001??: s4_gnt[7-1:0] = 7'b0000100;
   7'b000001?: s4_gnt[7-1:0] = 7'b0000010;
   7'b0000001: s4_gnt[7-1:0] = 7'b0000001;
   default: s4_gnt[7-1:0] = 7'b0000000;
endcase
end
assign s5_req_all[7-1:0] = s5_req[7-1:0] | s5_req_pend[7-1:0];
always @( s5_req_all[6:0])
begin
casez(s5_req_all[7-1:0])
   7'b1??????: s5_gnt[7-1:0] = 7'b1000000;
   7'b01?????: s5_gnt[7-1:0] = 7'b0100000;
   7'b001????: s5_gnt[7-1:0] = 7'b0010000;
   7'b0001???: s5_gnt[7-1:0] = 7'b0001000;
   7'b00001??: s5_gnt[7-1:0] = 7'b0000100;
   7'b000001?: s5_gnt[7-1:0] = 7'b0000010;
   7'b0000001: s5_gnt[7-1:0] = 7'b0000001;
   default: s5_gnt[7-1:0] = 7'b0000000;
endcase
end
assign s6_req_all[7-1:0] = s6_req[7-1:0] | s6_req_pend[7-1:0];
always @( s6_req_all[6:0])
begin
casez(s6_req_all[7-1:0])
   7'b1??????: s6_gnt[7-1:0] = 7'b1000000;
   7'b01?????: s6_gnt[7-1:0] = 7'b0100000;
   7'b001????: s6_gnt[7-1:0] = 7'b0010000;
   7'b0001???: s6_gnt[7-1:0] = 7'b0001000;
   7'b00001??: s6_gnt[7-1:0] = 7'b0000100;
   7'b000001?: s6_gnt[7-1:0] = 7'b0000010;
   7'b0000001: s6_gnt[7-1:0] = 7'b0000001;
   default: s6_gnt[7-1:0] = 7'b0000000;
endcase
end
assign s7_req_all[7-1:0] = s7_req[7-1:0] | s7_req_pend[7-1:0];
always @( s7_req_all[6:0])
begin
casez(s7_req_all[7-1:0])
   7'b1??????: s7_gnt[7-1:0] = 7'b1000000;
   7'b01?????: s7_gnt[7-1:0] = 7'b0100000;
   7'b001????: s7_gnt[7-1:0] = 7'b0010000;
   7'b0001???: s7_gnt[7-1:0] = 7'b0001000;
   7'b00001??: s7_gnt[7-1:0] = 7'b0000100;
   7'b000001?: s7_gnt[7-1:0] = 7'b0000010;
   7'b0000001: s7_gnt[7-1:0] = 7'b0000001;
   default: s7_gnt[7-1:0] = 7'b0000000;
endcase
end
assign s8_req_all[7-1:0] = s8_req[7-1:0] | s8_req_pend[7-1:0];
always @( s8_req_all[6:0])
begin
casez(s8_req_all[7-1:0])
   7'b1??????: s8_gnt[7-1:0] = 7'b1000000;
   7'b01?????: s8_gnt[7-1:0] = 7'b0100000;
   7'b001????: s8_gnt[7-1:0] = 7'b0010000;
   7'b0001???: s8_gnt[7-1:0] = 7'b0001000;
   7'b00001??: s8_gnt[7-1:0] = 7'b0000100;
   7'b000001?: s8_gnt[7-1:0] = 7'b0000010;
   7'b0000001: s8_gnt[7-1:0] = 7'b0000001;
   default: s8_gnt[7-1:0] = 7'b0000000;
endcase
end
assign s9_req_all[7-1:0] = s9_req[7-1:0] | s9_req_pend[7-1:0];
always @( s9_req_all[6:0])
begin
casez(s9_req_all[7-1:0])
   7'b1??????: s9_gnt[7-1:0] = 7'b1000000;
   7'b01?????: s9_gnt[7-1:0] = 7'b0100000;
   7'b001????: s9_gnt[7-1:0] = 7'b0010000;
   7'b0001???: s9_gnt[7-1:0] = 7'b0001000;
   7'b00001??: s9_gnt[7-1:0] = 7'b0000100;
   7'b000001?: s9_gnt[7-1:0] = 7'b0000010;
   7'b0000001: s9_gnt[7-1:0] = 7'b0000001;
   default: s9_gnt[7-1:0] = 7'b0000000;
endcase
end
assign s10_req_all[7-1:0] = s10_req[7-1:0] | s10_req_pend[7-1:0];
always @( s10_req_all[6:0])
begin
casez(s10_req_all[7-1:0])
   7'b1??????: s10_gnt[7-1:0] = 7'b1000000;
   7'b01?????: s10_gnt[7-1:0] = 7'b0100000;
   7'b001????: s10_gnt[7-1:0] = 7'b0010000;
   7'b0001???: s10_gnt[7-1:0] = 7'b0001000;
   7'b00001??: s10_gnt[7-1:0] = 7'b0000100;
   7'b000001?: s10_gnt[7-1:0] = 7'b0000010;
   7'b0000001: s10_gnt[7-1:0] = 7'b0000001;
   default: s10_gnt[7-1:0] = 7'b0000000;
endcase
end
assign s11_req_all[7-1:0] = s11_req[7-1:0] | s11_req_pend[7-1:0];
always @( s11_req_all[6:0])
begin
casez(s11_req_all[7-1:0])
   7'b1??????: s11_gnt[7-1:0] = 7'b1000000;
   7'b01?????: s11_gnt[7-1:0] = 7'b0100000;
   7'b001????: s11_gnt[7-1:0] = 7'b0010000;
   7'b0001???: s11_gnt[7-1:0] = 7'b0001000;
   7'b00001??: s11_gnt[7-1:0] = 7'b0000100;
   7'b000001?: s11_gnt[7-1:0] = 7'b0000010;
   7'b0000001: s11_gnt[7-1:0] = 7'b0000001;
   default: s11_gnt[7-1:0] = 7'b0000000;
endcase
end
assign m0_s0_sel = s0_gnt[6];
assign m0_s0_wt_sel = s0_req_all[6] & ~s0_gnt[6];
assign m0_s1_sel = s1_gnt[6];
assign m0_s1_wt_sel = s1_req_all[6] & ~s1_gnt[6];
assign m0_s2_sel = s2_gnt[6];
assign m0_s2_wt_sel = s2_req_all[6] & ~s2_gnt[6];
assign m0_s3_sel = s3_gnt[6];
assign m0_s3_wt_sel = s3_req_all[6] & ~s3_gnt[6];
assign m0_s4_sel = s4_gnt[6];
assign m0_s4_wt_sel = s4_req_all[6] & ~s4_gnt[6];
assign m0_s5_sel = s5_gnt[6];
assign m0_s5_wt_sel = s5_req_all[6] & ~s5_gnt[6];
assign m0_s6_sel = s6_gnt[6];
assign m0_s6_wt_sel = s6_req_all[6] & ~s6_gnt[6];
assign m0_s7_sel = s7_gnt[6];
assign m0_s7_wt_sel = s7_req_all[6] & ~s7_gnt[6];
assign m0_s8_sel = s8_gnt[6];
assign m0_s8_wt_sel = s8_req_all[6] & ~s8_gnt[6];
assign m0_s9_sel = s9_gnt[6];
assign m0_s9_wt_sel = s9_req_all[6] & ~s9_gnt[6];
assign m0_s10_sel = s10_gnt[6];
assign m0_s10_wt_sel = s10_req_all[6] & ~s10_gnt[6];
assign m0_s11_sel = s11_gnt[6];
assign m0_s11_wt_sel = s11_req_all[6] & ~s11_gnt[6];
assign m1_s0_sel = s0_gnt[5];
assign m1_s0_wt_sel = s0_req_all[5] & ~s0_gnt[5];
assign m1_s1_sel = s1_gnt[5];
assign m1_s1_wt_sel = s1_req_all[5] & ~s1_gnt[5];
assign m1_s2_sel = s2_gnt[5];
assign m1_s2_wt_sel = s2_req_all[5] & ~s2_gnt[5];
assign m1_s3_sel = s3_gnt[5];
assign m1_s3_wt_sel = s3_req_all[5] & ~s3_gnt[5];
assign m1_s4_sel = s4_gnt[5];
assign m1_s4_wt_sel = s4_req_all[5] & ~s4_gnt[5];
assign m1_s5_sel = s5_gnt[5];
assign m1_s5_wt_sel = s5_req_all[5] & ~s5_gnt[5];
assign m1_s6_sel = s6_gnt[5];
assign m1_s6_wt_sel = s6_req_all[5] & ~s6_gnt[5];
assign m1_s7_sel = s7_gnt[5];
assign m1_s7_wt_sel = s7_req_all[5] & ~s7_gnt[5];
assign m1_s8_sel = s8_gnt[5];
assign m1_s8_wt_sel = s8_req_all[5] & ~s8_gnt[5];
assign m1_s9_sel = s9_gnt[5];
assign m1_s9_wt_sel = s9_req_all[5] & ~s9_gnt[5];
assign m1_s10_sel = s10_gnt[5];
assign m1_s10_wt_sel = s10_req_all[5] & ~s10_gnt[5];
assign m1_s11_sel = s11_gnt[5];
assign m1_s11_wt_sel = s11_req_all[5] & ~s11_gnt[5];
assign m2_s0_sel = s0_gnt[4];
assign m2_s0_wt_sel = s0_req_all[4] & ~s0_gnt[4];
assign m2_s1_sel = s1_gnt[4];
assign m2_s1_wt_sel = s1_req_all[4] & ~s1_gnt[4];
assign m2_s2_sel = s2_gnt[4];
assign m2_s2_wt_sel = s2_req_all[4] & ~s2_gnt[4];
assign m2_s3_sel = s3_gnt[4];
assign m2_s3_wt_sel = s3_req_all[4] & ~s3_gnt[4];
assign m2_s4_sel = s4_gnt[4];
assign m2_s4_wt_sel = s4_req_all[4] & ~s4_gnt[4];
assign m2_s5_sel = s5_gnt[4];
assign m2_s5_wt_sel = s5_req_all[4] & ~s5_gnt[4];
assign m2_s6_sel = s6_gnt[4];
assign m2_s6_wt_sel = s6_req_all[4] & ~s6_gnt[4];
assign m2_s7_sel = s7_gnt[4];
assign m2_s7_wt_sel = s7_req_all[4] & ~s7_gnt[4];
assign m2_s8_sel = s8_gnt[4];
assign m2_s8_wt_sel = s8_req_all[4] & ~s8_gnt[4];
assign m2_s9_sel = s9_gnt[4];
assign m2_s9_wt_sel = s9_req_all[4] & ~s9_gnt[4];
assign m2_s10_sel = s10_gnt[4];
assign m2_s10_wt_sel = s10_req_all[4] & ~s10_gnt[4];
assign m2_s11_sel = s11_gnt[4];
assign m2_s11_wt_sel = s11_req_all[4] & ~s11_gnt[4];
assign m3_s0_sel = s0_gnt[3];
assign m3_s0_wt_sel = s0_req_all[3] & ~s0_gnt[3];
assign m3_s1_sel = s1_gnt[3];
assign m3_s1_wt_sel = s1_req_all[3] & ~s1_gnt[3];
assign m3_s2_sel = s2_gnt[3];
assign m3_s2_wt_sel = s2_req_all[3] & ~s2_gnt[3];
assign m3_s3_sel = s3_gnt[3];
assign m3_s3_wt_sel = s3_req_all[3] & ~s3_gnt[3];
assign m3_s4_sel = s4_gnt[3];
assign m3_s4_wt_sel = s4_req_all[3] & ~s4_gnt[3];
assign m3_s5_sel = s5_gnt[3];
assign m3_s5_wt_sel = s5_req_all[3] & ~s5_gnt[3];
assign m3_s6_sel = s6_gnt[3];
assign m3_s6_wt_sel = s6_req_all[3] & ~s6_gnt[3];
assign m3_s7_sel = s7_gnt[3];
assign m3_s7_wt_sel = s7_req_all[3] & ~s7_gnt[3];
assign m3_s8_sel = s8_gnt[3];
assign m3_s8_wt_sel = s8_req_all[3] & ~s8_gnt[3];
assign m3_s9_sel = s9_gnt[3];
assign m3_s9_wt_sel = s9_req_all[3] & ~s9_gnt[3];
assign m3_s10_sel = s10_gnt[3];
assign m3_s10_wt_sel = s10_req_all[3] & ~s10_gnt[3];
assign m3_s11_sel = s11_gnt[3];
assign m3_s11_wt_sel = s11_req_all[3] & ~s11_gnt[3];
assign m4_s0_sel = s0_gnt[2];
assign m4_s0_wt_sel = s0_req_all[2] & ~s0_gnt[2];
assign m4_s1_sel = s1_gnt[2];
assign m4_s1_wt_sel = s1_req_all[2] & ~s1_gnt[2];
assign m4_s2_sel = s2_gnt[2];
assign m4_s2_wt_sel = s2_req_all[2] & ~s2_gnt[2];
assign m4_s3_sel = s3_gnt[2];
assign m4_s3_wt_sel = s3_req_all[2] & ~s3_gnt[2];
assign m4_s4_sel = s4_gnt[2];
assign m4_s4_wt_sel = s4_req_all[2] & ~s4_gnt[2];
assign m4_s5_sel = s5_gnt[2];
assign m4_s5_wt_sel = s5_req_all[2] & ~s5_gnt[2];
assign m4_s6_sel = s6_gnt[2];
assign m4_s6_wt_sel = s6_req_all[2] & ~s6_gnt[2];
assign m4_s7_sel = s7_gnt[2];
assign m4_s7_wt_sel = s7_req_all[2] & ~s7_gnt[2];
assign m4_s8_sel = s8_gnt[2];
assign m4_s8_wt_sel = s8_req_all[2] & ~s8_gnt[2];
assign m4_s9_sel = s9_gnt[2];
assign m4_s9_wt_sel = s9_req_all[2] & ~s9_gnt[2];
assign m4_s10_sel = s10_gnt[2];
assign m4_s10_wt_sel = s10_req_all[2] & ~s10_gnt[2];
assign m4_s11_sel = s11_gnt[2];
assign m4_s11_wt_sel = s11_req_all[2] & ~s11_gnt[2];
assign m5_s0_sel = s0_gnt[1];
assign m5_s0_wt_sel = s0_req_all[1] & ~s0_gnt[1];
assign m5_s1_sel = s1_gnt[1];
assign m5_s1_wt_sel = s1_req_all[1] & ~s1_gnt[1];
assign m5_s2_sel = s2_gnt[1];
assign m5_s2_wt_sel = s2_req_all[1] & ~s2_gnt[1];
assign m5_s3_sel = s3_gnt[1];
assign m5_s3_wt_sel = s3_req_all[1] & ~s3_gnt[1];
assign m5_s4_sel = s4_gnt[1];
assign m5_s4_wt_sel = s4_req_all[1] & ~s4_gnt[1];
assign m5_s5_sel = s5_gnt[1];
assign m5_s5_wt_sel = s5_req_all[1] & ~s5_gnt[1];
assign m5_s6_sel = s6_gnt[1];
assign m5_s6_wt_sel = s6_req_all[1] & ~s6_gnt[1];
assign m5_s7_sel = s7_gnt[1];
assign m5_s7_wt_sel = s7_req_all[1] & ~s7_gnt[1];
assign m5_s8_sel = s8_gnt[1];
assign m5_s8_wt_sel = s8_req_all[1] & ~s8_gnt[1];
assign m5_s9_sel = s9_gnt[1];
assign m5_s9_wt_sel = s9_req_all[1] & ~s9_gnt[1];
assign m5_s10_sel = s10_gnt[1];
assign m5_s10_wt_sel = s10_req_all[1] & ~s10_gnt[1];
assign m5_s11_sel = s11_gnt[1];
assign m5_s11_wt_sel = s11_req_all[1] & ~s11_gnt[1];
assign m6_s0_sel = s0_gnt[0];
assign m6_s0_wt_sel = s0_req_all[0] & ~s0_gnt[0];
assign m6_s1_sel = s1_gnt[0];
assign m6_s1_wt_sel = s1_req_all[0] & ~s1_gnt[0];
assign m6_s2_sel = s2_gnt[0];
assign m6_s2_wt_sel = s2_req_all[0] & ~s2_gnt[0];
assign m6_s3_sel = s3_gnt[0];
assign m6_s3_wt_sel = s3_req_all[0] & ~s3_gnt[0];
assign m6_s4_sel = s4_gnt[0];
assign m6_s4_wt_sel = s4_req_all[0] & ~s4_gnt[0];
assign m6_s5_sel = s5_gnt[0];
assign m6_s5_wt_sel = s5_req_all[0] & ~s5_gnt[0];
assign m6_s6_sel = s6_gnt[0];
assign m6_s6_wt_sel = s6_req_all[0] & ~s6_gnt[0];
assign m6_s7_sel = s7_gnt[0];
assign m6_s7_wt_sel = s7_req_all[0] & ~s7_gnt[0];
assign m6_s8_sel = s8_gnt[0];
assign m6_s8_wt_sel = s8_req_all[0] & ~s8_gnt[0];
assign m6_s9_sel = s9_gnt[0];
assign m6_s9_wt_sel = s9_req_all[0] & ~s9_gnt[0];
assign m6_s10_sel = s10_gnt[0];
assign m6_s10_wt_sel = s10_req_all[0] & ~s10_gnt[0];
assign m6_s11_sel = s11_gnt[0];
assign m6_s11_wt_sel = s11_req_all[0] & ~s11_gnt[0];
assign m0_s0_hld =
                       (|m1_cur_st[4:3]) ||
                       (|m2_cur_st[4:3]) ||
                       (|m3_cur_st[4:3]) ||
                       (|m4_cur_st[4:3]) ||
                       (|m5_cur_st[4:3]) ||
                       (|m6_cur_st[4:3]);
assign m0_s1_hld =
                       (|m1_cur_st[8:7]) ||
                       (|m2_cur_st[8:7]) ||
                       (|m3_cur_st[8:7]) ||
                       (|m4_cur_st[8:7]) ||
                       (|m5_cur_st[8:7]) ||
                       (|m6_cur_st[8:7]);
assign m0_s2_hld =
                       (|m1_cur_st[12:11]) ||
                       (|m2_cur_st[12:11]) ||
                       (|m3_cur_st[12:11]) ||
                       (|m4_cur_st[12:11]) ||
                       (|m5_cur_st[12:11]) ||
                       (|m6_cur_st[12:11]);
assign m0_s3_hld =
                       (|m1_cur_st[16:15]) ||
                       (|m2_cur_st[16:15]) ||
                       (|m3_cur_st[16:15]) ||
                       (|m4_cur_st[16:15]) ||
                       (|m5_cur_st[16:15]) ||
                       (|m6_cur_st[16:15]);
assign m0_s4_hld =
                       (|m1_cur_st[20:19]) ||
                       (|m2_cur_st[20:19]) ||
                       (|m3_cur_st[20:19]) ||
                       (|m4_cur_st[20:19]) ||
                       (|m5_cur_st[20:19]) ||
                       (|m6_cur_st[20:19]);
assign m0_s5_hld =
                       (|m1_cur_st[24:23]) ||
                       (|m2_cur_st[24:23]) ||
                       (|m3_cur_st[24:23]) ||
                       (|m4_cur_st[24:23]) ||
                       (|m5_cur_st[24:23]) ||
                       (|m6_cur_st[24:23]);
assign m0_s6_hld =
                       (|m1_cur_st[28:27]) ||
                       (|m2_cur_st[28:27]) ||
                       (|m3_cur_st[28:27]) ||
                       (|m4_cur_st[28:27]) ||
                       (|m5_cur_st[28:27]) ||
                       (|m6_cur_st[28:27]);
assign m0_s7_hld =
                       (|m1_cur_st[32:31]) ||
                       (|m2_cur_st[32:31]) ||
                       (|m3_cur_st[32:31]) ||
                       (|m4_cur_st[32:31]) ||
                       (|m5_cur_st[32:31]) ||
                       (|m6_cur_st[32:31]);
assign m0_s8_hld =
                       (|m1_cur_st[36:35]) ||
                       (|m2_cur_st[36:35]) ||
                       (|m3_cur_st[36:35]) ||
                       (|m4_cur_st[36:35]) ||
                       (|m5_cur_st[36:35]) ||
                       (|m6_cur_st[36:35]);
assign m0_s9_hld =
                       (|m1_cur_st[40:39]) ||
                       (|m2_cur_st[40:39]) ||
                       (|m3_cur_st[40:39]) ||
                       (|m4_cur_st[40:39]) ||
                       (|m5_cur_st[40:39]) ||
                       (|m6_cur_st[40:39]);
assign m0_s10_hld =
                       (|m1_cur_st[44:43]) ||
                       (|m2_cur_st[44:43]) ||
                       (|m3_cur_st[44:43]) ||
                       (|m4_cur_st[44:43]) ||
                       (|m5_cur_st[44:43]) ||
                       (|m6_cur_st[44:43]);
assign m0_s11_hld =
                       (|m1_cur_st[48:47]) ||
                       (|m2_cur_st[48:47]) ||
                       (|m3_cur_st[48:47]) ||
                       (|m4_cur_st[48:47]) ||
                       (|m5_cur_st[48:47]) ||
                       (|m6_cur_st[48:47]);
assign m1_s0_hld =
                       (|m0_cur_st[4:3]) ||
                       (|m2_cur_st[4:3]) ||
                       (|m3_cur_st[4:3]) ||
                       (|m4_cur_st[4:3]) ||
                       (|m5_cur_st[4:3]) ||
                       (|m6_cur_st[4:3]);
assign m1_s1_hld =
                       (|m0_cur_st[8:7]) ||
                       (|m2_cur_st[8:7]) ||
                       (|m3_cur_st[8:7]) ||
                       (|m4_cur_st[8:7]) ||
                       (|m5_cur_st[8:7]) ||
                       (|m6_cur_st[8:7]);
assign m1_s2_hld =
                       (|m0_cur_st[12:11]) ||
                       (|m2_cur_st[12:11]) ||
                       (|m3_cur_st[12:11]) ||
                       (|m4_cur_st[12:11]) ||
                       (|m5_cur_st[12:11]) ||
                       (|m6_cur_st[12:11]);
assign m1_s3_hld =
                       (|m0_cur_st[16:15]) ||
                       (|m2_cur_st[16:15]) ||
                       (|m3_cur_st[16:15]) ||
                       (|m4_cur_st[16:15]) ||
                       (|m5_cur_st[16:15]) ||
                       (|m6_cur_st[16:15]);
assign m1_s4_hld =
                       (|m0_cur_st[20:19]) ||
                       (|m2_cur_st[20:19]) ||
                       (|m3_cur_st[20:19]) ||
                       (|m4_cur_st[20:19]) ||
                       (|m5_cur_st[20:19]) ||
                       (|m6_cur_st[20:19]);
assign m1_s5_hld =
                       (|m0_cur_st[24:23]) ||
                       (|m2_cur_st[24:23]) ||
                       (|m3_cur_st[24:23]) ||
                       (|m4_cur_st[24:23]) ||
                       (|m5_cur_st[24:23]) ||
                       (|m6_cur_st[24:23]);
assign m1_s6_hld =
                       (|m0_cur_st[28:27]) ||
                       (|m2_cur_st[28:27]) ||
                       (|m3_cur_st[28:27]) ||
                       (|m4_cur_st[28:27]) ||
                       (|m5_cur_st[28:27]) ||
                       (|m6_cur_st[28:27]);
assign m1_s7_hld =
                       (|m0_cur_st[32:31]) ||
                       (|m2_cur_st[32:31]) ||
                       (|m3_cur_st[32:31]) ||
                       (|m4_cur_st[32:31]) ||
                       (|m5_cur_st[32:31]) ||
                       (|m6_cur_st[32:31]);
assign m1_s8_hld =
                       (|m0_cur_st[36:35]) ||
                       (|m2_cur_st[36:35]) ||
                       (|m3_cur_st[36:35]) ||
                       (|m4_cur_st[36:35]) ||
                       (|m5_cur_st[36:35]) ||
                       (|m6_cur_st[36:35]);
assign m1_s9_hld =
                       (|m0_cur_st[40:39]) ||
                       (|m2_cur_st[40:39]) ||
                       (|m3_cur_st[40:39]) ||
                       (|m4_cur_st[40:39]) ||
                       (|m5_cur_st[40:39]) ||
                       (|m6_cur_st[40:39]);
assign m1_s10_hld =
                       (|m0_cur_st[44:43]) ||
                       (|m2_cur_st[44:43]) ||
                       (|m3_cur_st[44:43]) ||
                       (|m4_cur_st[44:43]) ||
                       (|m5_cur_st[44:43]) ||
                       (|m6_cur_st[44:43]);
assign m1_s11_hld =
                       (|m0_cur_st[48:47]) ||
                       (|m2_cur_st[48:47]) ||
                       (|m3_cur_st[48:47]) ||
                       (|m4_cur_st[48:47]) ||
                       (|m5_cur_st[48:47]) ||
                       (|m6_cur_st[48:47]);
assign m2_s0_hld =
                       (|m0_cur_st[4:3]) ||
                       (|m1_cur_st[4:3]) ||
                       (|m3_cur_st[4:3]) ||
                       (|m4_cur_st[4:3]) ||
                       (|m5_cur_st[4:3]) ||
                       (|m6_cur_st[4:3]);
assign m2_s1_hld =
                       (|m0_cur_st[8:7]) ||
                       (|m1_cur_st[8:7]) ||
                       (|m3_cur_st[8:7]) ||
                       (|m4_cur_st[8:7]) ||
                       (|m5_cur_st[8:7]) ||
                       (|m6_cur_st[8:7]);
assign m2_s2_hld =
                       (|m0_cur_st[12:11]) ||
                       (|m1_cur_st[12:11]) ||
                       (|m3_cur_st[12:11]) ||
                       (|m4_cur_st[12:11]) ||
                       (|m5_cur_st[12:11]) ||
                       (|m6_cur_st[12:11]);
assign m2_s3_hld =
                       (|m0_cur_st[16:15]) ||
                       (|m1_cur_st[16:15]) ||
                       (|m3_cur_st[16:15]) ||
                       (|m4_cur_st[16:15]) ||
                       (|m5_cur_st[16:15]) ||
                       (|m6_cur_st[16:15]);
assign m2_s4_hld =
                       (|m0_cur_st[20:19]) ||
                       (|m1_cur_st[20:19]) ||
                       (|m3_cur_st[20:19]) ||
                       (|m4_cur_st[20:19]) ||
                       (|m5_cur_st[20:19]) ||
                       (|m6_cur_st[20:19]);
assign m2_s5_hld =
                       (|m0_cur_st[24:23]) ||
                       (|m1_cur_st[24:23]) ||
                       (|m3_cur_st[24:23]) ||
                       (|m4_cur_st[24:23]) ||
                       (|m5_cur_st[24:23]) ||
                       (|m6_cur_st[24:23]);
assign m2_s6_hld =
                       (|m0_cur_st[28:27]) ||
                       (|m1_cur_st[28:27]) ||
                       (|m3_cur_st[28:27]) ||
                       (|m4_cur_st[28:27]) ||
                       (|m5_cur_st[28:27]) ||
                       (|m6_cur_st[28:27]);
assign m2_s7_hld =
                       (|m0_cur_st[32:31]) ||
                       (|m1_cur_st[32:31]) ||
                       (|m3_cur_st[32:31]) ||
                       (|m4_cur_st[32:31]) ||
                       (|m5_cur_st[32:31]) ||
                       (|m6_cur_st[32:31]);
assign m2_s8_hld =
                       (|m0_cur_st[36:35]) ||
                       (|m1_cur_st[36:35]) ||
                       (|m3_cur_st[36:35]) ||
                       (|m4_cur_st[36:35]) ||
                       (|m5_cur_st[36:35]) ||
                       (|m6_cur_st[36:35]);
assign m2_s9_hld =
                       (|m0_cur_st[40:39]) ||
                       (|m1_cur_st[40:39]) ||
                       (|m3_cur_st[40:39]) ||
                       (|m4_cur_st[40:39]) ||
                       (|m5_cur_st[40:39]) ||
                       (|m6_cur_st[40:39]);
assign m2_s10_hld =
                       (|m0_cur_st[44:43]) ||
                       (|m1_cur_st[44:43]) ||
                       (|m3_cur_st[44:43]) ||
                       (|m4_cur_st[44:43]) ||
                       (|m5_cur_st[44:43]) ||
                       (|m6_cur_st[44:43]);
assign m2_s11_hld =
                       (|m0_cur_st[48:47]) ||
                       (|m1_cur_st[48:47]) ||
                       (|m3_cur_st[48:47]) ||
                       (|m4_cur_st[48:47]) ||
                       (|m5_cur_st[48:47]) ||
                       (|m6_cur_st[48:47]);
assign m3_s0_hld =
                       (|m0_cur_st[4:3]) ||
                       (|m1_cur_st[4:3]) ||
                       (|m2_cur_st[4:3]) ||
                       (|m4_cur_st[4:3]) ||
                       (|m5_cur_st[4:3]) ||
                       (|m6_cur_st[4:3]);
assign m3_s1_hld =
                       (|m0_cur_st[8:7]) ||
                       (|m1_cur_st[8:7]) ||
                       (|m2_cur_st[8:7]) ||
                       (|m4_cur_st[8:7]) ||
                       (|m5_cur_st[8:7]) ||
                       (|m6_cur_st[8:7]);
assign m3_s2_hld =
                       (|m0_cur_st[12:11]) ||
                       (|m1_cur_st[12:11]) ||
                       (|m2_cur_st[12:11]) ||
                       (|m4_cur_st[12:11]) ||
                       (|m5_cur_st[12:11]) ||
                       (|m6_cur_st[12:11]);
assign m3_s3_hld =
                       (|m0_cur_st[16:15]) ||
                       (|m1_cur_st[16:15]) ||
                       (|m2_cur_st[16:15]) ||
                       (|m4_cur_st[16:15]) ||
                       (|m5_cur_st[16:15]) ||
                       (|m6_cur_st[16:15]);
assign m3_s4_hld =
                       (|m0_cur_st[20:19]) ||
                       (|m1_cur_st[20:19]) ||
                       (|m2_cur_st[20:19]) ||
                       (|m4_cur_st[20:19]) ||
                       (|m5_cur_st[20:19]) ||
                       (|m6_cur_st[20:19]);
assign m3_s5_hld =
                       (|m0_cur_st[24:23]) ||
                       (|m1_cur_st[24:23]) ||
                       (|m2_cur_st[24:23]) ||
                       (|m4_cur_st[24:23]) ||
                       (|m5_cur_st[24:23]) ||
                       (|m6_cur_st[24:23]);
assign m3_s6_hld =
                       (|m0_cur_st[28:27]) ||
                       (|m1_cur_st[28:27]) ||
                       (|m2_cur_st[28:27]) ||
                       (|m4_cur_st[28:27]) ||
                       (|m5_cur_st[28:27]) ||
                       (|m6_cur_st[28:27]);
assign m3_s7_hld =
                       (|m0_cur_st[32:31]) ||
                       (|m1_cur_st[32:31]) ||
                       (|m2_cur_st[32:31]) ||
                       (|m4_cur_st[32:31]) ||
                       (|m5_cur_st[32:31]) ||
                       (|m6_cur_st[32:31]);
assign m3_s8_hld =
                       (|m0_cur_st[36:35]) ||
                       (|m1_cur_st[36:35]) ||
                       (|m2_cur_st[36:35]) ||
                       (|m4_cur_st[36:35]) ||
                       (|m5_cur_st[36:35]) ||
                       (|m6_cur_st[36:35]);
assign m3_s9_hld =
                       (|m0_cur_st[40:39]) ||
                       (|m1_cur_st[40:39]) ||
                       (|m2_cur_st[40:39]) ||
                       (|m4_cur_st[40:39]) ||
                       (|m5_cur_st[40:39]) ||
                       (|m6_cur_st[40:39]);
assign m3_s10_hld =
                       (|m0_cur_st[44:43]) ||
                       (|m1_cur_st[44:43]) ||
                       (|m2_cur_st[44:43]) ||
                       (|m4_cur_st[44:43]) ||
                       (|m5_cur_st[44:43]) ||
                       (|m6_cur_st[44:43]);
assign m3_s11_hld =
                       (|m0_cur_st[48:47]) ||
                       (|m1_cur_st[48:47]) ||
                       (|m2_cur_st[48:47]) ||
                       (|m4_cur_st[48:47]) ||
                       (|m5_cur_st[48:47]) ||
                       (|m6_cur_st[48:47]);
assign m4_s0_hld =
                       (|m0_cur_st[4:3]) ||
                       (|m1_cur_st[4:3]) ||
                       (|m2_cur_st[4:3]) ||
                       (|m3_cur_st[4:3]) ||
                       (|m5_cur_st[4:3]) ||
                       (|m6_cur_st[4:3]);
assign m4_s1_hld =
                       (|m0_cur_st[8:7]) ||
                       (|m1_cur_st[8:7]) ||
                       (|m2_cur_st[8:7]) ||
                       (|m3_cur_st[8:7]) ||
                       (|m5_cur_st[8:7]) ||
                       (|m6_cur_st[8:7]);
assign m4_s2_hld =
                       (|m0_cur_st[12:11]) ||
                       (|m1_cur_st[12:11]) ||
                       (|m2_cur_st[12:11]) ||
                       (|m3_cur_st[12:11]) ||
                       (|m5_cur_st[12:11]) ||
                       (|m6_cur_st[12:11]);
assign m4_s3_hld =
                       (|m0_cur_st[16:15]) ||
                       (|m1_cur_st[16:15]) ||
                       (|m2_cur_st[16:15]) ||
                       (|m3_cur_st[16:15]) ||
                       (|m5_cur_st[16:15]) ||
                       (|m6_cur_st[16:15]);
assign m4_s4_hld =
                       (|m0_cur_st[20:19]) ||
                       (|m1_cur_st[20:19]) ||
                       (|m2_cur_st[20:19]) ||
                       (|m3_cur_st[20:19]) ||
                       (|m5_cur_st[20:19]) ||
                       (|m6_cur_st[20:19]);
assign m4_s5_hld =
                       (|m0_cur_st[24:23]) ||
                       (|m1_cur_st[24:23]) ||
                       (|m2_cur_st[24:23]) ||
                       (|m3_cur_st[24:23]) ||
                       (|m5_cur_st[24:23]) ||
                       (|m6_cur_st[24:23]);
assign m4_s6_hld =
                       (|m0_cur_st[28:27]) ||
                       (|m1_cur_st[28:27]) ||
                       (|m2_cur_st[28:27]) ||
                       (|m3_cur_st[28:27]) ||
                       (|m5_cur_st[28:27]) ||
                       (|m6_cur_st[28:27]);
assign m4_s7_hld =
                       (|m0_cur_st[32:31]) ||
                       (|m1_cur_st[32:31]) ||
                       (|m2_cur_st[32:31]) ||
                       (|m3_cur_st[32:31]) ||
                       (|m5_cur_st[32:31]) ||
                       (|m6_cur_st[32:31]);
assign m4_s8_hld =
                       (|m0_cur_st[36:35]) ||
                       (|m1_cur_st[36:35]) ||
                       (|m2_cur_st[36:35]) ||
                       (|m3_cur_st[36:35]) ||
                       (|m5_cur_st[36:35]) ||
                       (|m6_cur_st[36:35]);
assign m4_s9_hld =
                       (|m0_cur_st[40:39]) ||
                       (|m1_cur_st[40:39]) ||
                       (|m2_cur_st[40:39]) ||
                       (|m3_cur_st[40:39]) ||
                       (|m5_cur_st[40:39]) ||
                       (|m6_cur_st[40:39]);
assign m4_s10_hld =
                       (|m0_cur_st[44:43]) ||
                       (|m1_cur_st[44:43]) ||
                       (|m2_cur_st[44:43]) ||
                       (|m3_cur_st[44:43]) ||
                       (|m5_cur_st[44:43]) ||
                       (|m6_cur_st[44:43]);
assign m4_s11_hld =
                       (|m0_cur_st[48:47]) ||
                       (|m1_cur_st[48:47]) ||
                       (|m2_cur_st[48:47]) ||
                       (|m3_cur_st[48:47]) ||
                       (|m5_cur_st[48:47]) ||
                       (|m6_cur_st[48:47]);
assign m5_s0_hld =
                       (|m0_cur_st[4:3]) ||
                       (|m1_cur_st[4:3]) ||
                       (|m2_cur_st[4:3]) ||
                       (|m3_cur_st[4:3]) ||
                       (|m4_cur_st[4:3]) ||
                       (|m6_cur_st[4:3]);
assign m5_s1_hld =
                       (|m0_cur_st[8:7]) ||
                       (|m1_cur_st[8:7]) ||
                       (|m2_cur_st[8:7]) ||
                       (|m3_cur_st[8:7]) ||
                       (|m4_cur_st[8:7]) ||
                       (|m6_cur_st[8:7]);
assign m5_s2_hld =
                       (|m0_cur_st[12:11]) ||
                       (|m1_cur_st[12:11]) ||
                       (|m2_cur_st[12:11]) ||
                       (|m3_cur_st[12:11]) ||
                       (|m4_cur_st[12:11]) ||
                       (|m6_cur_st[12:11]);
assign m5_s3_hld =
                       (|m0_cur_st[16:15]) ||
                       (|m1_cur_st[16:15]) ||
                       (|m2_cur_st[16:15]) ||
                       (|m3_cur_st[16:15]) ||
                       (|m4_cur_st[16:15]) ||
                       (|m6_cur_st[16:15]);
assign m5_s4_hld =
                       (|m0_cur_st[20:19]) ||
                       (|m1_cur_st[20:19]) ||
                       (|m2_cur_st[20:19]) ||
                       (|m3_cur_st[20:19]) ||
                       (|m4_cur_st[20:19]) ||
                       (|m6_cur_st[20:19]);
assign m5_s5_hld =
                       (|m0_cur_st[24:23]) ||
                       (|m1_cur_st[24:23]) ||
                       (|m2_cur_st[24:23]) ||
                       (|m3_cur_st[24:23]) ||
                       (|m4_cur_st[24:23]) ||
                       (|m6_cur_st[24:23]);
assign m5_s6_hld =
                       (|m0_cur_st[28:27]) ||
                       (|m1_cur_st[28:27]) ||
                       (|m2_cur_st[28:27]) ||
                       (|m3_cur_st[28:27]) ||
                       (|m4_cur_st[28:27]) ||
                       (|m6_cur_st[28:27]);
assign m5_s7_hld =
                       (|m0_cur_st[32:31]) ||
                       (|m1_cur_st[32:31]) ||
                       (|m2_cur_st[32:31]) ||
                       (|m3_cur_st[32:31]) ||
                       (|m4_cur_st[32:31]) ||
                       (|m6_cur_st[32:31]);
assign m5_s8_hld =
                       (|m0_cur_st[36:35]) ||
                       (|m1_cur_st[36:35]) ||
                       (|m2_cur_st[36:35]) ||
                       (|m3_cur_st[36:35]) ||
                       (|m4_cur_st[36:35]) ||
                       (|m6_cur_st[36:35]);
assign m5_s9_hld =
                       (|m0_cur_st[40:39]) ||
                       (|m1_cur_st[40:39]) ||
                       (|m2_cur_st[40:39]) ||
                       (|m3_cur_st[40:39]) ||
                       (|m4_cur_st[40:39]) ||
                       (|m6_cur_st[40:39]);
assign m5_s10_hld =
                       (|m0_cur_st[44:43]) ||
                       (|m1_cur_st[44:43]) ||
                       (|m2_cur_st[44:43]) ||
                       (|m3_cur_st[44:43]) ||
                       (|m4_cur_st[44:43]) ||
                       (|m6_cur_st[44:43]);
assign m5_s11_hld =
                       (|m0_cur_st[48:47]) ||
                       (|m1_cur_st[48:47]) ||
                       (|m2_cur_st[48:47]) ||
                       (|m3_cur_st[48:47]) ||
                       (|m4_cur_st[48:47]) ||
                       (|m6_cur_st[48:47]);
assign m6_s0_hld =
                       (|m0_cur_st[4:3]) ||
                       (|m1_cur_st[4:3]) ||
                       (|m2_cur_st[4:3]) ||
                       (|m3_cur_st[4:3]) ||
                       (|m4_cur_st[4:3]) ||
                       (|m5_cur_st[4:3]);
assign m6_s1_hld =
                       (|m0_cur_st[8:7]) ||
                       (|m1_cur_st[8:7]) ||
                       (|m2_cur_st[8:7]) ||
                       (|m3_cur_st[8:7]) ||
                       (|m4_cur_st[8:7]) ||
                       (|m5_cur_st[8:7]);
assign m6_s2_hld =
                       (|m0_cur_st[12:11]) ||
                       (|m1_cur_st[12:11]) ||
                       (|m2_cur_st[12:11]) ||
                       (|m3_cur_st[12:11]) ||
                       (|m4_cur_st[12:11]) ||
                       (|m5_cur_st[12:11]);
assign m6_s3_hld =
                       (|m0_cur_st[16:15]) ||
                       (|m1_cur_st[16:15]) ||
                       (|m2_cur_st[16:15]) ||
                       (|m3_cur_st[16:15]) ||
                       (|m4_cur_st[16:15]) ||
                       (|m5_cur_st[16:15]);
assign m6_s4_hld =
                       (|m0_cur_st[20:19]) ||
                       (|m1_cur_st[20:19]) ||
                       (|m2_cur_st[20:19]) ||
                       (|m3_cur_st[20:19]) ||
                       (|m4_cur_st[20:19]) ||
                       (|m5_cur_st[20:19]);
assign m6_s5_hld =
                       (|m0_cur_st[24:23]) ||
                       (|m1_cur_st[24:23]) ||
                       (|m2_cur_st[24:23]) ||
                       (|m3_cur_st[24:23]) ||
                       (|m4_cur_st[24:23]) ||
                       (|m5_cur_st[24:23]);
assign m6_s6_hld =
                       (|m0_cur_st[28:27]) ||
                       (|m1_cur_st[28:27]) ||
                       (|m2_cur_st[28:27]) ||
                       (|m3_cur_st[28:27]) ||
                       (|m4_cur_st[28:27]) ||
                       (|m5_cur_st[28:27]);
assign m6_s7_hld =
                       (|m0_cur_st[32:31]) ||
                       (|m1_cur_st[32:31]) ||
                       (|m2_cur_st[32:31]) ||
                       (|m3_cur_st[32:31]) ||
                       (|m4_cur_st[32:31]) ||
                       (|m5_cur_st[32:31]);
assign m6_s8_hld =
                       (|m0_cur_st[36:35]) ||
                       (|m1_cur_st[36:35]) ||
                       (|m2_cur_st[36:35]) ||
                       (|m3_cur_st[36:35]) ||
                       (|m4_cur_st[36:35]) ||
                       (|m5_cur_st[36:35]);
assign m6_s9_hld =
                       (|m0_cur_st[40:39]) ||
                       (|m1_cur_st[40:39]) ||
                       (|m2_cur_st[40:39]) ||
                       (|m3_cur_st[40:39]) ||
                       (|m4_cur_st[40:39]) ||
                       (|m5_cur_st[40:39]);
assign m6_s10_hld =
                       (|m0_cur_st[44:43]) ||
                       (|m1_cur_st[44:43]) ||
                       (|m2_cur_st[44:43]) ||
                       (|m3_cur_st[44:43]) ||
                       (|m4_cur_st[44:43]) ||
                       (|m5_cur_st[44:43]);
assign m6_s11_hld =
                       (|m0_cur_st[48:47]) ||
                       (|m1_cur_st[48:47]) ||
                       (|m2_cur_st[48:47]) ||
                       (|m3_cur_st[48:47]) ||
                       (|m4_cur_st[48:47]) ||
                       (|m5_cur_st[48:47]);
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
       m0_cur_st[48:0] <= S_IDLE;
    else
       m0_cur_st[48:0] <= m0_nxt_st[48:0];
  end
always @ (*)
begin
case(m0_cur_st[48:0])
  S_IDLE:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       case(1'b1)
         m0_s0_sel: begin
                          m0_nxt_st[48:0] = m0_s0_hld ? S_S0_WAIT : (s0_hready ? S_S0_DATA : S_S0_CMD);
                          m0_latch_cmd = m0_s0_hld ? 1'b1 : (s0_hready ? 1'b0 : 1'b1);
                          m0_s0_cmd_cur = m0_s0_hld ? 1'b0 : (s0_hready ? 1'b1 : 1'b0);
                        end
         m0_s0_wt_sel: begin
                             m0_nxt_st[48:0] = S_S0_GNT;
                             m0_latch_cmd = 1'b1;
                           end
         m0_s1_sel: begin
                          m0_nxt_st[48:0] = m0_s1_hld ? S_S1_WAIT : (s1_hready ? S_S1_DATA : S_S1_CMD);
                          m0_latch_cmd = m0_s1_hld ? 1'b1 : (s1_hready ? 1'b0 : 1'b1);
                          m0_s1_cmd_cur = m0_s1_hld ? 1'b0 : (s1_hready ? 1'b1 : 1'b0);
                        end
         m0_s1_wt_sel: begin
                             m0_nxt_st[48:0] = S_S1_GNT;
                             m0_latch_cmd = 1'b1;
                           end
         m0_s2_sel: begin
                          m0_nxt_st[48:0] = m0_s2_hld ? S_S2_WAIT : (s2_hready ? S_S2_DATA : S_S2_CMD);
                          m0_latch_cmd = m0_s2_hld ? 1'b1 : (s2_hready ? 1'b0 : 1'b1);
                          m0_s2_cmd_cur = m0_s2_hld ? 1'b0 : (s2_hready ? 1'b1 : 1'b0);
                        end
         m0_s2_wt_sel: begin
                             m0_nxt_st[48:0] = S_S2_GNT;
                             m0_latch_cmd = 1'b1;
                           end
         m0_s3_sel: begin
                          m0_nxt_st[48:0] = m0_s3_hld ? S_S3_WAIT : (s3_hready ? S_S3_DATA : S_S3_CMD);
                          m0_latch_cmd = m0_s3_hld ? 1'b1 : (s3_hready ? 1'b0 : 1'b1);
                          m0_s3_cmd_cur = m0_s3_hld ? 1'b0 : (s3_hready ? 1'b1 : 1'b0);
                        end
         m0_s3_wt_sel: begin
                             m0_nxt_st[48:0] = S_S3_GNT;
                             m0_latch_cmd = 1'b1;
                           end
         m0_s4_sel: begin
                          m0_nxt_st[48:0] = m0_s4_hld ? S_S4_WAIT : (s4_hready ? S_S4_DATA : S_S4_CMD);
                          m0_latch_cmd = m0_s4_hld ? 1'b1 : (s4_hready ? 1'b0 : 1'b1);
                          m0_s4_cmd_cur = m0_s4_hld ? 1'b0 : (s4_hready ? 1'b1 : 1'b0);
                        end
         m0_s4_wt_sel: begin
                             m0_nxt_st[48:0] = S_S4_GNT;
                             m0_latch_cmd = 1'b1;
                           end
         m0_s5_sel: begin
                          m0_nxt_st[48:0] = m0_s5_hld ? S_S5_WAIT : (s5_hready ? S_S5_DATA : S_S5_CMD);
                          m0_latch_cmd = m0_s5_hld ? 1'b1 : (s5_hready ? 1'b0 : 1'b1);
                          m0_s5_cmd_cur = m0_s5_hld ? 1'b0 : (s5_hready ? 1'b1 : 1'b0);
                        end
         m0_s5_wt_sel: begin
                             m0_nxt_st[48:0] = S_S5_GNT;
                             m0_latch_cmd = 1'b1;
                           end
         m0_s6_sel: begin
                          m0_nxt_st[48:0] = m0_s6_hld ? S_S6_WAIT : (s6_hready ? S_S6_DATA : S_S6_CMD);
                          m0_latch_cmd = m0_s6_hld ? 1'b1 : (s6_hready ? 1'b0 : 1'b1);
                          m0_s6_cmd_cur = m0_s6_hld ? 1'b0 : (s6_hready ? 1'b1 : 1'b0);
                        end
         m0_s6_wt_sel: begin
                             m0_nxt_st[48:0] = S_S6_GNT;
                             m0_latch_cmd = 1'b1;
                           end
         m0_s7_sel: begin
                          m0_nxt_st[48:0] = m0_s7_hld ? S_S7_WAIT : (s7_hready ? S_S7_DATA : S_S7_CMD);
                          m0_latch_cmd = m0_s7_hld ? 1'b1 : (s7_hready ? 1'b0 : 1'b1);
                          m0_s7_cmd_cur = m0_s7_hld ? 1'b0 : (s7_hready ? 1'b1 : 1'b0);
                        end
         m0_s7_wt_sel: begin
                             m0_nxt_st[48:0] = S_S7_GNT;
                             m0_latch_cmd = 1'b1;
                           end
         m0_s8_sel: begin
                          m0_nxt_st[48:0] = m0_s8_hld ? S_S8_WAIT : (s8_hready ? S_S8_DATA : S_S8_CMD);
                          m0_latch_cmd = m0_s8_hld ? 1'b1 : (s8_hready ? 1'b0 : 1'b1);
                          m0_s8_cmd_cur = m0_s8_hld ? 1'b0 : (s8_hready ? 1'b1 : 1'b0);
                        end
         m0_s8_wt_sel: begin
                             m0_nxt_st[48:0] = S_S8_GNT;
                             m0_latch_cmd = 1'b1;
                           end
         m0_s9_sel: begin
                          m0_nxt_st[48:0] = m0_s9_hld ? S_S9_WAIT : (s9_hready ? S_S9_DATA : S_S9_CMD);
                          m0_latch_cmd = m0_s9_hld ? 1'b1 : (s9_hready ? 1'b0 : 1'b1);
                          m0_s9_cmd_cur = m0_s9_hld ? 1'b0 : (s9_hready ? 1'b1 : 1'b0);
                        end
         m0_s9_wt_sel: begin
                             m0_nxt_st[48:0] = S_S9_GNT;
                             m0_latch_cmd = 1'b1;
                           end
         m0_s10_sel: begin
                          m0_nxt_st[48:0] = m0_s10_hld ? S_S10_WAIT : (s10_hready ? S_S10_DATA : S_S10_CMD);
                          m0_latch_cmd = m0_s10_hld ? 1'b1 : (s10_hready ? 1'b0 : 1'b1);
                          m0_s10_cmd_cur = m0_s10_hld ? 1'b0 : (s10_hready ? 1'b1 : 1'b0);
                        end
         m0_s10_wt_sel: begin
                             m0_nxt_st[48:0] = S_S10_GNT;
                             m0_latch_cmd = 1'b1;
                           end
         m0_s11_sel: begin
                          m0_nxt_st[48:0] = m0_s11_hld ? S_S11_WAIT : (s11_hready ? S_S11_DATA : S_S11_CMD);
                          m0_latch_cmd = m0_s11_hld ? 1'b1 : (s11_hready ? 1'b0 : 1'b1);
                          m0_s11_cmd_cur = m0_s11_hld ? 1'b0 : (s11_hready ? 1'b1 : 1'b0);
                        end
         m0_s11_wt_sel: begin
                             m0_nxt_st[48:0] = S_S11_GNT;
                             m0_latch_cmd = 1'b1;
                           end
         default: begin
                          m0_nxt_st[48:0] = S_IDLE;
                  end
       endcase
  end
  S_S0_GNT:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       case(1'b1)
         m0_s0_sel: begin
                          m0_nxt_st[48:0] = m0_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                          m0_s0_cmd_last = m0_s0_hld ? 1'b0 : (s0_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m0_nxt_st[48:0] = S_S0_GNT;
                  end
       endcase
  end
  S_S1_GNT:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       case(1'b1)
         m0_s1_sel: begin
                          m0_nxt_st[48:0] = m0_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                          m0_s1_cmd_last = m0_s1_hld ? 1'b0 : (s1_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m0_nxt_st[48:0] = S_S1_GNT;
                  end
       endcase
  end
  S_S2_GNT:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       case(1'b1)
         m0_s2_sel: begin
                          m0_nxt_st[48:0] = m0_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                          m0_s2_cmd_last = m0_s2_hld ? 1'b0 : (s2_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m0_nxt_st[48:0] = S_S2_GNT;
                  end
       endcase
  end
  S_S3_GNT:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       case(1'b1)
         m0_s3_sel: begin
                          m0_nxt_st[48:0] = m0_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                          m0_s3_cmd_last = m0_s3_hld ? 1'b0 : (s3_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m0_nxt_st[48:0] = S_S3_GNT;
                  end
       endcase
  end
  S_S4_GNT:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       case(1'b1)
         m0_s4_sel: begin
                          m0_nxt_st[48:0] = m0_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                          m0_s4_cmd_last = m0_s4_hld ? 1'b0 : (s4_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m0_nxt_st[48:0] = S_S4_GNT;
                  end
       endcase
  end
  S_S5_GNT:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       case(1'b1)
         m0_s5_sel: begin
                          m0_nxt_st[48:0] = m0_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                          m0_s5_cmd_last = m0_s5_hld ? 1'b0 : (s5_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m0_nxt_st[48:0] = S_S5_GNT;
                  end
       endcase
  end
  S_S6_GNT:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       case(1'b1)
         m0_s6_sel: begin
                          m0_nxt_st[48:0] = m0_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                          m0_s6_cmd_last = m0_s6_hld ? 1'b0 : (s6_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m0_nxt_st[48:0] = S_S6_GNT;
                  end
       endcase
  end
  S_S7_GNT:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       case(1'b1)
         m0_s7_sel: begin
                          m0_nxt_st[48:0] = m0_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                          m0_s7_cmd_last = m0_s7_hld ? 1'b0 : (s7_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m0_nxt_st[48:0] = S_S7_GNT;
                  end
       endcase
  end
  S_S8_GNT:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       case(1'b1)
         m0_s8_sel: begin
                          m0_nxt_st[48:0] = m0_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                          m0_s8_cmd_last = m0_s8_hld ? 1'b0 : (s8_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m0_nxt_st[48:0] = S_S8_GNT;
                  end
       endcase
  end
  S_S9_GNT:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       case(1'b1)
         m0_s9_sel: begin
                          m0_nxt_st[48:0] = m0_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                          m0_s9_cmd_last = m0_s9_hld ? 1'b0 : (s9_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m0_nxt_st[48:0] = S_S9_GNT;
                  end
       endcase
  end
  S_S10_GNT:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       case(1'b1)
         m0_s10_sel: begin
                          m0_nxt_st[48:0] = m0_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                          m0_s10_cmd_last = m0_s10_hld ? 1'b0 : (s10_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m0_nxt_st[48:0] = S_S10_GNT;
                  end
       endcase
  end
  S_S11_GNT:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       case(1'b1)
         m0_s11_sel: begin
                          m0_nxt_st[48:0] = m0_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                          m0_s11_cmd_last = m0_s11_hld ? 1'b0 : (s11_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m0_nxt_st[48:0] = S_S11_GNT;
                  end
       endcase
  end
  S_S0_WAIT:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       case(1'b1)
         ~m0_s0_hld: begin
                          m0_nxt_st[48:0] = m0_s0_wt_sel ? S_S0_GNT : s0_hready ? S_S0_DATA : S_S0_CMD;
                          m0_s0_cmd_last = m0_s0_wt_sel ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m0_nxt_st[48:0] = S_S0_WAIT;
                  end
       endcase
  end
  S_S1_WAIT:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       case(1'b1)
         ~m0_s1_hld: begin
                          m0_nxt_st[48:0] = m0_s1_wt_sel ? S_S1_GNT : s1_hready ? S_S1_DATA : S_S1_CMD;
                          m0_s1_cmd_last = m0_s1_wt_sel ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m0_nxt_st[48:0] = S_S1_WAIT;
                  end
       endcase
  end
  S_S2_WAIT:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       case(1'b1)
         ~m0_s2_hld: begin
                          m0_nxt_st[48:0] = m0_s2_wt_sel ? S_S2_GNT : s2_hready ? S_S2_DATA : S_S2_CMD;
                          m0_s2_cmd_last = m0_s2_wt_sel ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m0_nxt_st[48:0] = S_S2_WAIT;
                  end
       endcase
  end
  S_S3_WAIT:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       case(1'b1)
         ~m0_s3_hld: begin
                          m0_nxt_st[48:0] = m0_s3_wt_sel ? S_S3_GNT : s3_hready ? S_S3_DATA : S_S3_CMD;
                          m0_s3_cmd_last = m0_s3_wt_sel ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m0_nxt_st[48:0] = S_S3_WAIT;
                  end
       endcase
  end
  S_S4_WAIT:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       case(1'b1)
         ~m0_s4_hld: begin
                          m0_nxt_st[48:0] = m0_s4_wt_sel ? S_S4_GNT : s4_hready ? S_S4_DATA : S_S4_CMD;
                          m0_s4_cmd_last = m0_s4_wt_sel ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m0_nxt_st[48:0] = S_S4_WAIT;
                  end
       endcase
  end
  S_S5_WAIT:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       case(1'b1)
         ~m0_s5_hld: begin
                          m0_nxt_st[48:0] = m0_s5_wt_sel ? S_S5_GNT : s5_hready ? S_S5_DATA : S_S5_CMD;
                          m0_s5_cmd_last = m0_s5_wt_sel ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m0_nxt_st[48:0] = S_S5_WAIT;
                  end
       endcase
  end
  S_S6_WAIT:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       case(1'b1)
         ~m0_s6_hld: begin
                          m0_nxt_st[48:0] = m0_s6_wt_sel ? S_S6_GNT : s6_hready ? S_S6_DATA : S_S6_CMD;
                          m0_s6_cmd_last = m0_s6_wt_sel ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m0_nxt_st[48:0] = S_S6_WAIT;
                  end
       endcase
  end
  S_S7_WAIT:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       case(1'b1)
         ~m0_s7_hld: begin
                          m0_nxt_st[48:0] = m0_s7_wt_sel ? S_S7_GNT : s7_hready ? S_S7_DATA : S_S7_CMD;
                          m0_s7_cmd_last = m0_s7_wt_sel ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m0_nxt_st[48:0] = S_S7_WAIT;
                  end
       endcase
  end
  S_S8_WAIT:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       case(1'b1)
         ~m0_s8_hld: begin
                          m0_nxt_st[48:0] = m0_s8_wt_sel ? S_S8_GNT : s8_hready ? S_S8_DATA : S_S8_CMD;
                          m0_s8_cmd_last = m0_s8_wt_sel ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m0_nxt_st[48:0] = S_S8_WAIT;
                  end
       endcase
  end
  S_S9_WAIT:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       case(1'b1)
         ~m0_s9_hld: begin
                          m0_nxt_st[48:0] = m0_s9_wt_sel ? S_S9_GNT : s9_hready ? S_S9_DATA : S_S9_CMD;
                          m0_s9_cmd_last = m0_s9_wt_sel ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m0_nxt_st[48:0] = S_S9_WAIT;
                  end
       endcase
  end
  S_S10_WAIT:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       case(1'b1)
         ~m0_s10_hld: begin
                          m0_nxt_st[48:0] = m0_s10_wt_sel ? S_S10_GNT : s10_hready ? S_S10_DATA : S_S10_CMD;
                          m0_s10_cmd_last = m0_s10_wt_sel ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m0_nxt_st[48:0] = S_S10_WAIT;
                  end
       endcase
  end
  S_S11_WAIT:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       case(1'b1)
         ~m0_s11_hld: begin
                          m0_nxt_st[48:0] = m0_s11_wt_sel ? S_S11_GNT : s11_hready ? S_S11_DATA : S_S11_CMD;
                          m0_s11_cmd_last = m0_s11_wt_sel ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m0_nxt_st[48:0] = S_S11_WAIT;
                  end
       endcase
  end
  S_S0_CMD: begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = s0_hready ? 1'b1 : 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       m0_nxt_st[48:0] = s0_hready  ? S_S0_DATA : S_S0_CMD;
  end
  S_S0_DATA:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b1;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       if(s0_hready)
         begin
           case(1'b1)
             m0_s0_sel: begin
                              m0_nxt_st[48:0] = S_S0_DATA;
                              m0_s0_cmd_cur = 1'b1;
                             end
             m0_s0_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S0_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s1_sel: begin
                              m0_nxt_st[48:0] = m0_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m0_latch_cmd = m0_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m0_s1_cmd_cur = m0_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m0_s1_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S1_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s2_sel: begin
                              m0_nxt_st[48:0] = m0_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m0_latch_cmd = m0_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m0_s2_cmd_cur = m0_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m0_s2_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S2_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s3_sel: begin
                              m0_nxt_st[48:0] = m0_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m0_latch_cmd = m0_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m0_s3_cmd_cur = m0_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m0_s3_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S3_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s4_sel: begin
                              m0_nxt_st[48:0] = m0_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m0_latch_cmd = m0_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m0_s4_cmd_cur = m0_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m0_s4_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S4_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s5_sel: begin
                              m0_nxt_st[48:0] = m0_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m0_latch_cmd = m0_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m0_s5_cmd_cur = m0_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m0_s5_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S5_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s6_sel: begin
                              m0_nxt_st[48:0] = m0_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m0_latch_cmd = m0_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m0_s6_cmd_cur = m0_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m0_s6_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S6_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s7_sel: begin
                              m0_nxt_st[48:0] = m0_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m0_latch_cmd = m0_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m0_s7_cmd_cur = m0_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m0_s7_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S7_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s8_sel: begin
                              m0_nxt_st[48:0] = m0_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m0_latch_cmd = m0_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m0_s8_cmd_cur = m0_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m0_s8_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S8_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s9_sel: begin
                              m0_nxt_st[48:0] = m0_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m0_latch_cmd = m0_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m0_s9_cmd_cur = m0_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m0_s9_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S9_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s10_sel: begin
                              m0_nxt_st[48:0] = m0_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m0_latch_cmd = m0_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m0_s10_cmd_cur = m0_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m0_s10_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S10_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s11_sel: begin
                              m0_nxt_st[48:0] = m0_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m0_latch_cmd = m0_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m0_s11_cmd_cur = m0_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m0_s11_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S11_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             default: begin
                             m0_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m0_nxt_st[48:0] = S_S0_DATA;
end
  S_S1_CMD: begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = s1_hready ? 1'b1 : 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       m0_nxt_st[48:0] = s1_hready  ? S_S1_DATA : S_S1_CMD;
  end
  S_S1_DATA:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b1;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       if(s1_hready)
         begin
           case(1'b1)
             m0_s0_sel: begin
                              m0_nxt_st[48:0] = m0_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m0_latch_cmd = m0_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m0_s0_cmd_cur = m0_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m0_s0_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S0_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s1_sel: begin
                              m0_nxt_st[48:0] = S_S1_DATA;
                              m0_s1_cmd_cur = 1'b1;
                             end
             m0_s1_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S1_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s2_sel: begin
                              m0_nxt_st[48:0] = m0_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m0_latch_cmd = m0_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m0_s2_cmd_cur = m0_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m0_s2_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S2_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s3_sel: begin
                              m0_nxt_st[48:0] = m0_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m0_latch_cmd = m0_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m0_s3_cmd_cur = m0_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m0_s3_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S3_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s4_sel: begin
                              m0_nxt_st[48:0] = m0_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m0_latch_cmd = m0_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m0_s4_cmd_cur = m0_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m0_s4_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S4_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s5_sel: begin
                              m0_nxt_st[48:0] = m0_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m0_latch_cmd = m0_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m0_s5_cmd_cur = m0_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m0_s5_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S5_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s6_sel: begin
                              m0_nxt_st[48:0] = m0_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m0_latch_cmd = m0_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m0_s6_cmd_cur = m0_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m0_s6_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S6_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s7_sel: begin
                              m0_nxt_st[48:0] = m0_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m0_latch_cmd = m0_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m0_s7_cmd_cur = m0_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m0_s7_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S7_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s8_sel: begin
                              m0_nxt_st[48:0] = m0_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m0_latch_cmd = m0_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m0_s8_cmd_cur = m0_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m0_s8_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S8_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s9_sel: begin
                              m0_nxt_st[48:0] = m0_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m0_latch_cmd = m0_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m0_s9_cmd_cur = m0_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m0_s9_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S9_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s10_sel: begin
                              m0_nxt_st[48:0] = m0_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m0_latch_cmd = m0_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m0_s10_cmd_cur = m0_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m0_s10_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S10_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s11_sel: begin
                              m0_nxt_st[48:0] = m0_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m0_latch_cmd = m0_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m0_s11_cmd_cur = m0_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m0_s11_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S11_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             default: begin
                             m0_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m0_nxt_st[48:0] = S_S1_DATA;
end
  S_S2_CMD: begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = s2_hready ? 1'b1 : 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       m0_nxt_st[48:0] = s2_hready  ? S_S2_DATA : S_S2_CMD;
  end
  S_S2_DATA:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b1;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       if(s2_hready)
         begin
           case(1'b1)
             m0_s0_sel: begin
                              m0_nxt_st[48:0] = m0_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m0_latch_cmd = m0_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m0_s0_cmd_cur = m0_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m0_s0_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S0_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s1_sel: begin
                              m0_nxt_st[48:0] = m0_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m0_latch_cmd = m0_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m0_s1_cmd_cur = m0_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m0_s1_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S1_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s2_sel: begin
                              m0_nxt_st[48:0] = S_S2_DATA;
                              m0_s2_cmd_cur = 1'b1;
                             end
             m0_s2_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S2_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s3_sel: begin
                              m0_nxt_st[48:0] = m0_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m0_latch_cmd = m0_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m0_s3_cmd_cur = m0_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m0_s3_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S3_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s4_sel: begin
                              m0_nxt_st[48:0] = m0_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m0_latch_cmd = m0_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m0_s4_cmd_cur = m0_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m0_s4_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S4_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s5_sel: begin
                              m0_nxt_st[48:0] = m0_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m0_latch_cmd = m0_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m0_s5_cmd_cur = m0_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m0_s5_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S5_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s6_sel: begin
                              m0_nxt_st[48:0] = m0_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m0_latch_cmd = m0_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m0_s6_cmd_cur = m0_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m0_s6_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S6_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s7_sel: begin
                              m0_nxt_st[48:0] = m0_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m0_latch_cmd = m0_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m0_s7_cmd_cur = m0_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m0_s7_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S7_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s8_sel: begin
                              m0_nxt_st[48:0] = m0_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m0_latch_cmd = m0_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m0_s8_cmd_cur = m0_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m0_s8_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S8_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s9_sel: begin
                              m0_nxt_st[48:0] = m0_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m0_latch_cmd = m0_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m0_s9_cmd_cur = m0_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m0_s9_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S9_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s10_sel: begin
                              m0_nxt_st[48:0] = m0_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m0_latch_cmd = m0_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m0_s10_cmd_cur = m0_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m0_s10_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S10_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s11_sel: begin
                              m0_nxt_st[48:0] = m0_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m0_latch_cmd = m0_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m0_s11_cmd_cur = m0_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m0_s11_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S11_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             default: begin
                             m0_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m0_nxt_st[48:0] = S_S2_DATA;
end
  S_S3_CMD: begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = s3_hready ? 1'b1 : 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       m0_nxt_st[48:0] = s3_hready  ? S_S3_DATA : S_S3_CMD;
  end
  S_S3_DATA:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b1;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       if(s3_hready)
         begin
           case(1'b1)
             m0_s0_sel: begin
                              m0_nxt_st[48:0] = m0_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m0_latch_cmd = m0_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m0_s0_cmd_cur = m0_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m0_s0_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S0_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s1_sel: begin
                              m0_nxt_st[48:0] = m0_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m0_latch_cmd = m0_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m0_s1_cmd_cur = m0_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m0_s1_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S1_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s2_sel: begin
                              m0_nxt_st[48:0] = m0_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m0_latch_cmd = m0_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m0_s2_cmd_cur = m0_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m0_s2_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S2_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s3_sel: begin
                              m0_nxt_st[48:0] = S_S3_DATA;
                              m0_s3_cmd_cur = 1'b1;
                             end
             m0_s3_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S3_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s4_sel: begin
                              m0_nxt_st[48:0] = m0_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m0_latch_cmd = m0_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m0_s4_cmd_cur = m0_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m0_s4_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S4_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s5_sel: begin
                              m0_nxt_st[48:0] = m0_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m0_latch_cmd = m0_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m0_s5_cmd_cur = m0_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m0_s5_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S5_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s6_sel: begin
                              m0_nxt_st[48:0] = m0_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m0_latch_cmd = m0_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m0_s6_cmd_cur = m0_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m0_s6_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S6_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s7_sel: begin
                              m0_nxt_st[48:0] = m0_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m0_latch_cmd = m0_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m0_s7_cmd_cur = m0_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m0_s7_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S7_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s8_sel: begin
                              m0_nxt_st[48:0] = m0_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m0_latch_cmd = m0_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m0_s8_cmd_cur = m0_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m0_s8_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S8_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s9_sel: begin
                              m0_nxt_st[48:0] = m0_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m0_latch_cmd = m0_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m0_s9_cmd_cur = m0_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m0_s9_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S9_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s10_sel: begin
                              m0_nxt_st[48:0] = m0_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m0_latch_cmd = m0_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m0_s10_cmd_cur = m0_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m0_s10_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S10_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s11_sel: begin
                              m0_nxt_st[48:0] = m0_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m0_latch_cmd = m0_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m0_s11_cmd_cur = m0_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m0_s11_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S11_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             default: begin
                             m0_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m0_nxt_st[48:0] = S_S3_DATA;
end
  S_S4_CMD: begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = s4_hready ? 1'b1 : 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       m0_nxt_st[48:0] = s4_hready  ? S_S4_DATA : S_S4_CMD;
  end
  S_S4_DATA:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b1;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       if(s4_hready)
         begin
           case(1'b1)
             m0_s0_sel: begin
                              m0_nxt_st[48:0] = m0_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m0_latch_cmd = m0_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m0_s0_cmd_cur = m0_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m0_s0_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S0_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s1_sel: begin
                              m0_nxt_st[48:0] = m0_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m0_latch_cmd = m0_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m0_s1_cmd_cur = m0_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m0_s1_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S1_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s2_sel: begin
                              m0_nxt_st[48:0] = m0_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m0_latch_cmd = m0_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m0_s2_cmd_cur = m0_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m0_s2_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S2_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s3_sel: begin
                              m0_nxt_st[48:0] = m0_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m0_latch_cmd = m0_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m0_s3_cmd_cur = m0_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m0_s3_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S3_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s4_sel: begin
                              m0_nxt_st[48:0] = S_S4_DATA;
                              m0_s4_cmd_cur = 1'b1;
                             end
             m0_s4_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S4_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s5_sel: begin
                              m0_nxt_st[48:0] = m0_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m0_latch_cmd = m0_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m0_s5_cmd_cur = m0_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m0_s5_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S5_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s6_sel: begin
                              m0_nxt_st[48:0] = m0_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m0_latch_cmd = m0_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m0_s6_cmd_cur = m0_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m0_s6_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S6_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s7_sel: begin
                              m0_nxt_st[48:0] = m0_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m0_latch_cmd = m0_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m0_s7_cmd_cur = m0_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m0_s7_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S7_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s8_sel: begin
                              m0_nxt_st[48:0] = m0_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m0_latch_cmd = m0_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m0_s8_cmd_cur = m0_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m0_s8_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S8_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s9_sel: begin
                              m0_nxt_st[48:0] = m0_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m0_latch_cmd = m0_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m0_s9_cmd_cur = m0_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m0_s9_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S9_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s10_sel: begin
                              m0_nxt_st[48:0] = m0_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m0_latch_cmd = m0_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m0_s10_cmd_cur = m0_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m0_s10_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S10_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s11_sel: begin
                              m0_nxt_st[48:0] = m0_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m0_latch_cmd = m0_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m0_s11_cmd_cur = m0_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m0_s11_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S11_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             default: begin
                             m0_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m0_nxt_st[48:0] = S_S4_DATA;
end
  S_S5_CMD: begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = s5_hready ? 1'b1 : 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       m0_nxt_st[48:0] = s5_hready  ? S_S5_DATA : S_S5_CMD;
  end
  S_S5_DATA:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b1;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       if(s5_hready)
         begin
           case(1'b1)
             m0_s0_sel: begin
                              m0_nxt_st[48:0] = m0_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m0_latch_cmd = m0_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m0_s0_cmd_cur = m0_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m0_s0_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S0_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s1_sel: begin
                              m0_nxt_st[48:0] = m0_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m0_latch_cmd = m0_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m0_s1_cmd_cur = m0_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m0_s1_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S1_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s2_sel: begin
                              m0_nxt_st[48:0] = m0_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m0_latch_cmd = m0_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m0_s2_cmd_cur = m0_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m0_s2_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S2_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s3_sel: begin
                              m0_nxt_st[48:0] = m0_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m0_latch_cmd = m0_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m0_s3_cmd_cur = m0_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m0_s3_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S3_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s4_sel: begin
                              m0_nxt_st[48:0] = m0_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m0_latch_cmd = m0_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m0_s4_cmd_cur = m0_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m0_s4_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S4_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s5_sel: begin
                              m0_nxt_st[48:0] = S_S5_DATA;
                              m0_s5_cmd_cur = 1'b1;
                             end
             m0_s5_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S5_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s6_sel: begin
                              m0_nxt_st[48:0] = m0_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m0_latch_cmd = m0_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m0_s6_cmd_cur = m0_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m0_s6_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S6_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s7_sel: begin
                              m0_nxt_st[48:0] = m0_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m0_latch_cmd = m0_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m0_s7_cmd_cur = m0_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m0_s7_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S7_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s8_sel: begin
                              m0_nxt_st[48:0] = m0_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m0_latch_cmd = m0_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m0_s8_cmd_cur = m0_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m0_s8_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S8_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s9_sel: begin
                              m0_nxt_st[48:0] = m0_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m0_latch_cmd = m0_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m0_s9_cmd_cur = m0_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m0_s9_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S9_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s10_sel: begin
                              m0_nxt_st[48:0] = m0_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m0_latch_cmd = m0_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m0_s10_cmd_cur = m0_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m0_s10_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S10_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s11_sel: begin
                              m0_nxt_st[48:0] = m0_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m0_latch_cmd = m0_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m0_s11_cmd_cur = m0_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m0_s11_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S11_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             default: begin
                             m0_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m0_nxt_st[48:0] = S_S5_DATA;
end
  S_S6_CMD: begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = s6_hready ? 1'b1 : 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       m0_nxt_st[48:0] = s6_hready  ? S_S6_DATA : S_S6_CMD;
  end
  S_S6_DATA:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b1;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       if(s6_hready)
         begin
           case(1'b1)
             m0_s0_sel: begin
                              m0_nxt_st[48:0] = m0_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m0_latch_cmd = m0_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m0_s0_cmd_cur = m0_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m0_s0_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S0_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s1_sel: begin
                              m0_nxt_st[48:0] = m0_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m0_latch_cmd = m0_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m0_s1_cmd_cur = m0_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m0_s1_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S1_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s2_sel: begin
                              m0_nxt_st[48:0] = m0_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m0_latch_cmd = m0_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m0_s2_cmd_cur = m0_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m0_s2_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S2_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s3_sel: begin
                              m0_nxt_st[48:0] = m0_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m0_latch_cmd = m0_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m0_s3_cmd_cur = m0_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m0_s3_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S3_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s4_sel: begin
                              m0_nxt_st[48:0] = m0_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m0_latch_cmd = m0_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m0_s4_cmd_cur = m0_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m0_s4_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S4_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s5_sel: begin
                              m0_nxt_st[48:0] = m0_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m0_latch_cmd = m0_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m0_s5_cmd_cur = m0_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m0_s5_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S5_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s6_sel: begin
                              m0_nxt_st[48:0] = S_S6_DATA;
                              m0_s6_cmd_cur = 1'b1;
                             end
             m0_s6_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S6_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s7_sel: begin
                              m0_nxt_st[48:0] = m0_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m0_latch_cmd = m0_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m0_s7_cmd_cur = m0_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m0_s7_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S7_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s8_sel: begin
                              m0_nxt_st[48:0] = m0_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m0_latch_cmd = m0_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m0_s8_cmd_cur = m0_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m0_s8_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S8_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s9_sel: begin
                              m0_nxt_st[48:0] = m0_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m0_latch_cmd = m0_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m0_s9_cmd_cur = m0_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m0_s9_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S9_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s10_sel: begin
                              m0_nxt_st[48:0] = m0_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m0_latch_cmd = m0_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m0_s10_cmd_cur = m0_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m0_s10_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S10_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s11_sel: begin
                              m0_nxt_st[48:0] = m0_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m0_latch_cmd = m0_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m0_s11_cmd_cur = m0_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m0_s11_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S11_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             default: begin
                             m0_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m0_nxt_st[48:0] = S_S6_DATA;
end
  S_S7_CMD: begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = s7_hready ? 1'b1 : 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       m0_nxt_st[48:0] = s7_hready  ? S_S7_DATA : S_S7_CMD;
  end
  S_S7_DATA:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b1;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       if(s7_hready)
         begin
           case(1'b1)
             m0_s0_sel: begin
                              m0_nxt_st[48:0] = m0_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m0_latch_cmd = m0_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m0_s0_cmd_cur = m0_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m0_s0_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S0_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s1_sel: begin
                              m0_nxt_st[48:0] = m0_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m0_latch_cmd = m0_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m0_s1_cmd_cur = m0_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m0_s1_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S1_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s2_sel: begin
                              m0_nxt_st[48:0] = m0_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m0_latch_cmd = m0_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m0_s2_cmd_cur = m0_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m0_s2_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S2_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s3_sel: begin
                              m0_nxt_st[48:0] = m0_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m0_latch_cmd = m0_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m0_s3_cmd_cur = m0_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m0_s3_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S3_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s4_sel: begin
                              m0_nxt_st[48:0] = m0_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m0_latch_cmd = m0_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m0_s4_cmd_cur = m0_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m0_s4_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S4_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s5_sel: begin
                              m0_nxt_st[48:0] = m0_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m0_latch_cmd = m0_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m0_s5_cmd_cur = m0_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m0_s5_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S5_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s6_sel: begin
                              m0_nxt_st[48:0] = m0_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m0_latch_cmd = m0_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m0_s6_cmd_cur = m0_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m0_s6_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S6_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s7_sel: begin
                              m0_nxt_st[48:0] = S_S7_DATA;
                              m0_s7_cmd_cur = 1'b1;
                             end
             m0_s7_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S7_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s8_sel: begin
                              m0_nxt_st[48:0] = m0_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m0_latch_cmd = m0_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m0_s8_cmd_cur = m0_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m0_s8_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S8_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s9_sel: begin
                              m0_nxt_st[48:0] = m0_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m0_latch_cmd = m0_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m0_s9_cmd_cur = m0_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m0_s9_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S9_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s10_sel: begin
                              m0_nxt_st[48:0] = m0_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m0_latch_cmd = m0_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m0_s10_cmd_cur = m0_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m0_s10_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S10_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s11_sel: begin
                              m0_nxt_st[48:0] = m0_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m0_latch_cmd = m0_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m0_s11_cmd_cur = m0_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m0_s11_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S11_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             default: begin
                             m0_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m0_nxt_st[48:0] = S_S7_DATA;
end
  S_S8_CMD: begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = s8_hready ? 1'b1 : 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       m0_nxt_st[48:0] = s8_hready  ? S_S8_DATA : S_S8_CMD;
  end
  S_S8_DATA:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b1;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       if(s8_hready)
         begin
           case(1'b1)
             m0_s0_sel: begin
                              m0_nxt_st[48:0] = m0_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m0_latch_cmd = m0_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m0_s0_cmd_cur = m0_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m0_s0_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S0_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s1_sel: begin
                              m0_nxt_st[48:0] = m0_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m0_latch_cmd = m0_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m0_s1_cmd_cur = m0_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m0_s1_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S1_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s2_sel: begin
                              m0_nxt_st[48:0] = m0_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m0_latch_cmd = m0_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m0_s2_cmd_cur = m0_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m0_s2_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S2_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s3_sel: begin
                              m0_nxt_st[48:0] = m0_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m0_latch_cmd = m0_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m0_s3_cmd_cur = m0_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m0_s3_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S3_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s4_sel: begin
                              m0_nxt_st[48:0] = m0_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m0_latch_cmd = m0_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m0_s4_cmd_cur = m0_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m0_s4_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S4_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s5_sel: begin
                              m0_nxt_st[48:0] = m0_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m0_latch_cmd = m0_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m0_s5_cmd_cur = m0_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m0_s5_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S5_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s6_sel: begin
                              m0_nxt_st[48:0] = m0_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m0_latch_cmd = m0_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m0_s6_cmd_cur = m0_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m0_s6_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S6_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s7_sel: begin
                              m0_nxt_st[48:0] = m0_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m0_latch_cmd = m0_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m0_s7_cmd_cur = m0_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m0_s7_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S7_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s8_sel: begin
                              m0_nxt_st[48:0] = S_S8_DATA;
                              m0_s8_cmd_cur = 1'b1;
                             end
             m0_s8_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S8_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s9_sel: begin
                              m0_nxt_st[48:0] = m0_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m0_latch_cmd = m0_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m0_s9_cmd_cur = m0_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m0_s9_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S9_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s10_sel: begin
                              m0_nxt_st[48:0] = m0_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m0_latch_cmd = m0_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m0_s10_cmd_cur = m0_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m0_s10_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S10_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s11_sel: begin
                              m0_nxt_st[48:0] = m0_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m0_latch_cmd = m0_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m0_s11_cmd_cur = m0_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m0_s11_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S11_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             default: begin
                             m0_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m0_nxt_st[48:0] = S_S8_DATA;
end
  S_S9_CMD: begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = s9_hready ? 1'b1 : 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       m0_nxt_st[48:0] = s9_hready  ? S_S9_DATA : S_S9_CMD;
  end
  S_S9_DATA:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b1;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       if(s9_hready)
         begin
           case(1'b1)
             m0_s0_sel: begin
                              m0_nxt_st[48:0] = m0_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m0_latch_cmd = m0_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m0_s0_cmd_cur = m0_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m0_s0_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S0_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s1_sel: begin
                              m0_nxt_st[48:0] = m0_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m0_latch_cmd = m0_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m0_s1_cmd_cur = m0_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m0_s1_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S1_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s2_sel: begin
                              m0_nxt_st[48:0] = m0_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m0_latch_cmd = m0_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m0_s2_cmd_cur = m0_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m0_s2_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S2_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s3_sel: begin
                              m0_nxt_st[48:0] = m0_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m0_latch_cmd = m0_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m0_s3_cmd_cur = m0_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m0_s3_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S3_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s4_sel: begin
                              m0_nxt_st[48:0] = m0_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m0_latch_cmd = m0_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m0_s4_cmd_cur = m0_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m0_s4_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S4_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s5_sel: begin
                              m0_nxt_st[48:0] = m0_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m0_latch_cmd = m0_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m0_s5_cmd_cur = m0_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m0_s5_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S5_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s6_sel: begin
                              m0_nxt_st[48:0] = m0_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m0_latch_cmd = m0_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m0_s6_cmd_cur = m0_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m0_s6_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S6_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s7_sel: begin
                              m0_nxt_st[48:0] = m0_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m0_latch_cmd = m0_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m0_s7_cmd_cur = m0_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m0_s7_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S7_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s8_sel: begin
                              m0_nxt_st[48:0] = m0_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m0_latch_cmd = m0_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m0_s8_cmd_cur = m0_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m0_s8_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S8_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s9_sel: begin
                              m0_nxt_st[48:0] = S_S9_DATA;
                              m0_s9_cmd_cur = 1'b1;
                             end
             m0_s9_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S9_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s10_sel: begin
                              m0_nxt_st[48:0] = m0_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m0_latch_cmd = m0_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m0_s10_cmd_cur = m0_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m0_s10_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S10_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s11_sel: begin
                              m0_nxt_st[48:0] = m0_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m0_latch_cmd = m0_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m0_s11_cmd_cur = m0_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m0_s11_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S11_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             default: begin
                             m0_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m0_nxt_st[48:0] = S_S9_DATA;
end
  S_S10_CMD: begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = s10_hready ? 1'b1 : 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       m0_nxt_st[48:0] = s10_hready  ? S_S10_DATA : S_S10_CMD;
  end
  S_S10_DATA:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b1;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       if(s10_hready)
         begin
           case(1'b1)
             m0_s0_sel: begin
                              m0_nxt_st[48:0] = m0_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m0_latch_cmd = m0_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m0_s0_cmd_cur = m0_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m0_s0_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S0_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s1_sel: begin
                              m0_nxt_st[48:0] = m0_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m0_latch_cmd = m0_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m0_s1_cmd_cur = m0_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m0_s1_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S1_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s2_sel: begin
                              m0_nxt_st[48:0] = m0_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m0_latch_cmd = m0_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m0_s2_cmd_cur = m0_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m0_s2_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S2_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s3_sel: begin
                              m0_nxt_st[48:0] = m0_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m0_latch_cmd = m0_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m0_s3_cmd_cur = m0_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m0_s3_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S3_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s4_sel: begin
                              m0_nxt_st[48:0] = m0_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m0_latch_cmd = m0_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m0_s4_cmd_cur = m0_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m0_s4_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S4_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s5_sel: begin
                              m0_nxt_st[48:0] = m0_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m0_latch_cmd = m0_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m0_s5_cmd_cur = m0_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m0_s5_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S5_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s6_sel: begin
                              m0_nxt_st[48:0] = m0_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m0_latch_cmd = m0_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m0_s6_cmd_cur = m0_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m0_s6_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S6_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s7_sel: begin
                              m0_nxt_st[48:0] = m0_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m0_latch_cmd = m0_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m0_s7_cmd_cur = m0_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m0_s7_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S7_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s8_sel: begin
                              m0_nxt_st[48:0] = m0_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m0_latch_cmd = m0_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m0_s8_cmd_cur = m0_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m0_s8_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S8_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s9_sel: begin
                              m0_nxt_st[48:0] = m0_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m0_latch_cmd = m0_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m0_s9_cmd_cur = m0_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m0_s9_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S9_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s10_sel: begin
                              m0_nxt_st[48:0] = S_S10_DATA;
                              m0_s10_cmd_cur = 1'b1;
                             end
             m0_s10_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S10_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s11_sel: begin
                              m0_nxt_st[48:0] = m0_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m0_latch_cmd = m0_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m0_s11_cmd_cur = m0_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m0_s11_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S11_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             default: begin
                             m0_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m0_nxt_st[48:0] = S_S10_DATA;
end
  S_S11_CMD: begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = s11_hready ? 1'b1 : 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b0;
       m0_nxt_st[48:0] = s11_hready  ? S_S11_DATA : S_S11_CMD;
  end
  S_S11_DATA:begin
       m0_latch_cmd = 1'b0;
       m0_s0_cmd_last = 1'b0;
       m0_s0_cmd_cur = 1'b0;
       m0_s0_data = 1'b0;
       m0_s1_cmd_last = 1'b0;
       m0_s1_cmd_cur = 1'b0;
       m0_s1_data = 1'b0;
       m0_s2_cmd_last = 1'b0;
       m0_s2_cmd_cur = 1'b0;
       m0_s2_data = 1'b0;
       m0_s3_cmd_last = 1'b0;
       m0_s3_cmd_cur = 1'b0;
       m0_s3_data = 1'b0;
       m0_s4_cmd_last = 1'b0;
       m0_s4_cmd_cur = 1'b0;
       m0_s4_data = 1'b0;
       m0_s5_cmd_last = 1'b0;
       m0_s5_cmd_cur = 1'b0;
       m0_s5_data = 1'b0;
       m0_s6_cmd_last = 1'b0;
       m0_s6_cmd_cur = 1'b0;
       m0_s6_data = 1'b0;
       m0_s7_cmd_last = 1'b0;
       m0_s7_cmd_cur = 1'b0;
       m0_s7_data = 1'b0;
       m0_s8_cmd_last = 1'b0;
       m0_s8_cmd_cur = 1'b0;
       m0_s8_data = 1'b0;
       m0_s9_cmd_last = 1'b0;
       m0_s9_cmd_cur = 1'b0;
       m0_s9_data = 1'b0;
       m0_s10_cmd_last = 1'b0;
       m0_s10_cmd_cur = 1'b0;
       m0_s10_data = 1'b0;
       m0_s11_cmd_last = 1'b0;
       m0_s11_cmd_cur = 1'b0;
       m0_s11_data = 1'b1;
       if(s11_hready)
         begin
           case(1'b1)
             m0_s0_sel: begin
                              m0_nxt_st[48:0] = m0_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m0_latch_cmd = m0_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m0_s0_cmd_cur = m0_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m0_s0_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S0_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s1_sel: begin
                              m0_nxt_st[48:0] = m0_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m0_latch_cmd = m0_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m0_s1_cmd_cur = m0_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m0_s1_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S1_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s2_sel: begin
                              m0_nxt_st[48:0] = m0_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m0_latch_cmd = m0_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m0_s2_cmd_cur = m0_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m0_s2_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S2_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s3_sel: begin
                              m0_nxt_st[48:0] = m0_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m0_latch_cmd = m0_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m0_s3_cmd_cur = m0_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m0_s3_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S3_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s4_sel: begin
                              m0_nxt_st[48:0] = m0_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m0_latch_cmd = m0_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m0_s4_cmd_cur = m0_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m0_s4_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S4_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s5_sel: begin
                              m0_nxt_st[48:0] = m0_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m0_latch_cmd = m0_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m0_s5_cmd_cur = m0_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m0_s5_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S5_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s6_sel: begin
                              m0_nxt_st[48:0] = m0_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m0_latch_cmd = m0_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m0_s6_cmd_cur = m0_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m0_s6_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S6_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s7_sel: begin
                              m0_nxt_st[48:0] = m0_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m0_latch_cmd = m0_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m0_s7_cmd_cur = m0_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m0_s7_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S7_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s8_sel: begin
                              m0_nxt_st[48:0] = m0_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m0_latch_cmd = m0_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m0_s8_cmd_cur = m0_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m0_s8_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S8_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s9_sel: begin
                              m0_nxt_st[48:0] = m0_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m0_latch_cmd = m0_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m0_s9_cmd_cur = m0_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m0_s9_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S9_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s10_sel: begin
                              m0_nxt_st[48:0] = m0_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m0_latch_cmd = m0_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m0_s10_cmd_cur = m0_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m0_s10_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S10_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             m0_s11_sel: begin
                              m0_nxt_st[48:0] = S_S11_DATA;
                              m0_s11_cmd_cur = 1'b1;
                             end
             m0_s11_wt_sel: begin
                                 m0_nxt_st[48:0] = S_S11_GNT;
                                 m0_latch_cmd = 1'b1;
                               end
             default: begin
                             m0_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m0_nxt_st[48:0] = S_S11_DATA;
end
  default: begin
             m0_latch_cmd = 1'b0;
             m0_s0_cmd_last = 1'b0;
             m0_s0_cmd_cur = 1'b0;
             m0_s0_data = 1'b0;
             m0_s1_cmd_last = 1'b0;
             m0_s1_cmd_cur = 1'b0;
             m0_s1_data = 1'b0;
             m0_s2_cmd_last = 1'b0;
             m0_s2_cmd_cur = 1'b0;
             m0_s2_data = 1'b0;
             m0_s3_cmd_last = 1'b0;
             m0_s3_cmd_cur = 1'b0;
             m0_s3_data = 1'b0;
             m0_s4_cmd_last = 1'b0;
             m0_s4_cmd_cur = 1'b0;
             m0_s4_data = 1'b0;
             m0_s5_cmd_last = 1'b0;
             m0_s5_cmd_cur = 1'b0;
             m0_s5_data = 1'b0;
             m0_s6_cmd_last = 1'b0;
             m0_s6_cmd_cur = 1'b0;
             m0_s6_data = 1'b0;
             m0_s7_cmd_last = 1'b0;
             m0_s7_cmd_cur = 1'b0;
             m0_s7_data = 1'b0;
             m0_s8_cmd_last = 1'b0;
             m0_s8_cmd_cur = 1'b0;
             m0_s8_data = 1'b0;
             m0_s9_cmd_last = 1'b0;
             m0_s9_cmd_cur = 1'b0;
             m0_s9_data = 1'b0;
             m0_s10_cmd_last = 1'b0;
             m0_s10_cmd_cur = 1'b0;
             m0_s10_data = 1'b0;
             m0_s11_cmd_last = 1'b0;
             m0_s11_cmd_cur = 1'b0;
             m0_s11_data = 1'b0;
             m0_nxt_st[48:0] = S_IDLE;
  end
endcase
end
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
       m1_cur_st[48:0] <= S_IDLE;
    else
       m1_cur_st[48:0] <= m1_nxt_st[48:0];
  end
always @ (*)
begin
case(m1_cur_st[48:0])
  S_IDLE:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       case(1'b1)
         m1_s0_sel: begin
                          m1_nxt_st[48:0] = m1_s0_hld ? S_S0_WAIT : (s0_hready ? S_S0_DATA : S_S0_CMD);
                          m1_latch_cmd = m1_s0_hld ? 1'b1 : (s0_hready ? 1'b0 : 1'b1);
                          m1_s0_cmd_cur = m1_s0_hld ? 1'b0 : (s0_hready ? 1'b1 : 1'b0);
                        end
         m1_s0_wt_sel: begin
                             m1_nxt_st[48:0] = S_S0_GNT;
                             m1_latch_cmd = 1'b1;
                           end
         m1_s1_sel: begin
                          m1_nxt_st[48:0] = m1_s1_hld ? S_S1_WAIT : (s1_hready ? S_S1_DATA : S_S1_CMD);
                          m1_latch_cmd = m1_s1_hld ? 1'b1 : (s1_hready ? 1'b0 : 1'b1);
                          m1_s1_cmd_cur = m1_s1_hld ? 1'b0 : (s1_hready ? 1'b1 : 1'b0);
                        end
         m1_s1_wt_sel: begin
                             m1_nxt_st[48:0] = S_S1_GNT;
                             m1_latch_cmd = 1'b1;
                           end
         m1_s2_sel: begin
                          m1_nxt_st[48:0] = m1_s2_hld ? S_S2_WAIT : (s2_hready ? S_S2_DATA : S_S2_CMD);
                          m1_latch_cmd = m1_s2_hld ? 1'b1 : (s2_hready ? 1'b0 : 1'b1);
                          m1_s2_cmd_cur = m1_s2_hld ? 1'b0 : (s2_hready ? 1'b1 : 1'b0);
                        end
         m1_s2_wt_sel: begin
                             m1_nxt_st[48:0] = S_S2_GNT;
                             m1_latch_cmd = 1'b1;
                           end
         m1_s3_sel: begin
                          m1_nxt_st[48:0] = m1_s3_hld ? S_S3_WAIT : (s3_hready ? S_S3_DATA : S_S3_CMD);
                          m1_latch_cmd = m1_s3_hld ? 1'b1 : (s3_hready ? 1'b0 : 1'b1);
                          m1_s3_cmd_cur = m1_s3_hld ? 1'b0 : (s3_hready ? 1'b1 : 1'b0);
                        end
         m1_s3_wt_sel: begin
                             m1_nxt_st[48:0] = S_S3_GNT;
                             m1_latch_cmd = 1'b1;
                           end
         m1_s4_sel: begin
                          m1_nxt_st[48:0] = m1_s4_hld ? S_S4_WAIT : (s4_hready ? S_S4_DATA : S_S4_CMD);
                          m1_latch_cmd = m1_s4_hld ? 1'b1 : (s4_hready ? 1'b0 : 1'b1);
                          m1_s4_cmd_cur = m1_s4_hld ? 1'b0 : (s4_hready ? 1'b1 : 1'b0);
                        end
         m1_s4_wt_sel: begin
                             m1_nxt_st[48:0] = S_S4_GNT;
                             m1_latch_cmd = 1'b1;
                           end
         m1_s5_sel: begin
                          m1_nxt_st[48:0] = m1_s5_hld ? S_S5_WAIT : (s5_hready ? S_S5_DATA : S_S5_CMD);
                          m1_latch_cmd = m1_s5_hld ? 1'b1 : (s5_hready ? 1'b0 : 1'b1);
                          m1_s5_cmd_cur = m1_s5_hld ? 1'b0 : (s5_hready ? 1'b1 : 1'b0);
                        end
         m1_s5_wt_sel: begin
                             m1_nxt_st[48:0] = S_S5_GNT;
                             m1_latch_cmd = 1'b1;
                           end
         m1_s6_sel: begin
                          m1_nxt_st[48:0] = m1_s6_hld ? S_S6_WAIT : (s6_hready ? S_S6_DATA : S_S6_CMD);
                          m1_latch_cmd = m1_s6_hld ? 1'b1 : (s6_hready ? 1'b0 : 1'b1);
                          m1_s6_cmd_cur = m1_s6_hld ? 1'b0 : (s6_hready ? 1'b1 : 1'b0);
                        end
         m1_s6_wt_sel: begin
                             m1_nxt_st[48:0] = S_S6_GNT;
                             m1_latch_cmd = 1'b1;
                           end
         m1_s7_sel: begin
                          m1_nxt_st[48:0] = m1_s7_hld ? S_S7_WAIT : (s7_hready ? S_S7_DATA : S_S7_CMD);
                          m1_latch_cmd = m1_s7_hld ? 1'b1 : (s7_hready ? 1'b0 : 1'b1);
                          m1_s7_cmd_cur = m1_s7_hld ? 1'b0 : (s7_hready ? 1'b1 : 1'b0);
                        end
         m1_s7_wt_sel: begin
                             m1_nxt_st[48:0] = S_S7_GNT;
                             m1_latch_cmd = 1'b1;
                           end
         m1_s8_sel: begin
                          m1_nxt_st[48:0] = m1_s8_hld ? S_S8_WAIT : (s8_hready ? S_S8_DATA : S_S8_CMD);
                          m1_latch_cmd = m1_s8_hld ? 1'b1 : (s8_hready ? 1'b0 : 1'b1);
                          m1_s8_cmd_cur = m1_s8_hld ? 1'b0 : (s8_hready ? 1'b1 : 1'b0);
                        end
         m1_s8_wt_sel: begin
                             m1_nxt_st[48:0] = S_S8_GNT;
                             m1_latch_cmd = 1'b1;
                           end
         m1_s9_sel: begin
                          m1_nxt_st[48:0] = m1_s9_hld ? S_S9_WAIT : (s9_hready ? S_S9_DATA : S_S9_CMD);
                          m1_latch_cmd = m1_s9_hld ? 1'b1 : (s9_hready ? 1'b0 : 1'b1);
                          m1_s9_cmd_cur = m1_s9_hld ? 1'b0 : (s9_hready ? 1'b1 : 1'b0);
                        end
         m1_s9_wt_sel: begin
                             m1_nxt_st[48:0] = S_S9_GNT;
                             m1_latch_cmd = 1'b1;
                           end
         m1_s10_sel: begin
                          m1_nxt_st[48:0] = m1_s10_hld ? S_S10_WAIT : (s10_hready ? S_S10_DATA : S_S10_CMD);
                          m1_latch_cmd = m1_s10_hld ? 1'b1 : (s10_hready ? 1'b0 : 1'b1);
                          m1_s10_cmd_cur = m1_s10_hld ? 1'b0 : (s10_hready ? 1'b1 : 1'b0);
                        end
         m1_s10_wt_sel: begin
                             m1_nxt_st[48:0] = S_S10_GNT;
                             m1_latch_cmd = 1'b1;
                           end
         m1_s11_sel: begin
                          m1_nxt_st[48:0] = m1_s11_hld ? S_S11_WAIT : (s11_hready ? S_S11_DATA : S_S11_CMD);
                          m1_latch_cmd = m1_s11_hld ? 1'b1 : (s11_hready ? 1'b0 : 1'b1);
                          m1_s11_cmd_cur = m1_s11_hld ? 1'b0 : (s11_hready ? 1'b1 : 1'b0);
                        end
         m1_s11_wt_sel: begin
                             m1_nxt_st[48:0] = S_S11_GNT;
                             m1_latch_cmd = 1'b1;
                           end
         default: begin
                          m1_nxt_st[48:0] = S_IDLE;
                  end
       endcase
  end
  S_S0_GNT:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       case(1'b1)
         m1_s0_sel: begin
                          m1_nxt_st[48:0] = m1_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                          m1_s0_cmd_last = m1_s0_hld ? 1'b0 : (s0_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m1_nxt_st[48:0] = S_S0_GNT;
                  end
       endcase
  end
  S_S1_GNT:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       case(1'b1)
         m1_s1_sel: begin
                          m1_nxt_st[48:0] = m1_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                          m1_s1_cmd_last = m1_s1_hld ? 1'b0 : (s1_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m1_nxt_st[48:0] = S_S1_GNT;
                  end
       endcase
  end
  S_S2_GNT:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       case(1'b1)
         m1_s2_sel: begin
                          m1_nxt_st[48:0] = m1_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                          m1_s2_cmd_last = m1_s2_hld ? 1'b0 : (s2_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m1_nxt_st[48:0] = S_S2_GNT;
                  end
       endcase
  end
  S_S3_GNT:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       case(1'b1)
         m1_s3_sel: begin
                          m1_nxt_st[48:0] = m1_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                          m1_s3_cmd_last = m1_s3_hld ? 1'b0 : (s3_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m1_nxt_st[48:0] = S_S3_GNT;
                  end
       endcase
  end
  S_S4_GNT:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       case(1'b1)
         m1_s4_sel: begin
                          m1_nxt_st[48:0] = m1_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                          m1_s4_cmd_last = m1_s4_hld ? 1'b0 : (s4_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m1_nxt_st[48:0] = S_S4_GNT;
                  end
       endcase
  end
  S_S5_GNT:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       case(1'b1)
         m1_s5_sel: begin
                          m1_nxt_st[48:0] = m1_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                          m1_s5_cmd_last = m1_s5_hld ? 1'b0 : (s5_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m1_nxt_st[48:0] = S_S5_GNT;
                  end
       endcase
  end
  S_S6_GNT:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       case(1'b1)
         m1_s6_sel: begin
                          m1_nxt_st[48:0] = m1_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                          m1_s6_cmd_last = m1_s6_hld ? 1'b0 : (s6_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m1_nxt_st[48:0] = S_S6_GNT;
                  end
       endcase
  end
  S_S7_GNT:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       case(1'b1)
         m1_s7_sel: begin
                          m1_nxt_st[48:0] = m1_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                          m1_s7_cmd_last = m1_s7_hld ? 1'b0 : (s7_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m1_nxt_st[48:0] = S_S7_GNT;
                  end
       endcase
  end
  S_S8_GNT:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       case(1'b1)
         m1_s8_sel: begin
                          m1_nxt_st[48:0] = m1_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                          m1_s8_cmd_last = m1_s8_hld ? 1'b0 : (s8_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m1_nxt_st[48:0] = S_S8_GNT;
                  end
       endcase
  end
  S_S9_GNT:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       case(1'b1)
         m1_s9_sel: begin
                          m1_nxt_st[48:0] = m1_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                          m1_s9_cmd_last = m1_s9_hld ? 1'b0 : (s9_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m1_nxt_st[48:0] = S_S9_GNT;
                  end
       endcase
  end
  S_S10_GNT:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       case(1'b1)
         m1_s10_sel: begin
                          m1_nxt_st[48:0] = m1_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                          m1_s10_cmd_last = m1_s10_hld ? 1'b0 : (s10_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m1_nxt_st[48:0] = S_S10_GNT;
                  end
       endcase
  end
  S_S11_GNT:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       case(1'b1)
         m1_s11_sel: begin
                          m1_nxt_st[48:0] = m1_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                          m1_s11_cmd_last = m1_s11_hld ? 1'b0 : (s11_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m1_nxt_st[48:0] = S_S11_GNT;
                  end
       endcase
  end
  S_S0_WAIT:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       case(1'b1)
         ~m1_s0_hld: begin
                          m1_nxt_st[48:0] = m1_s0_wt_sel ? S_S0_GNT : s0_hready ? S_S0_DATA : S_S0_CMD;
                          m1_s0_cmd_last = m1_s0_wt_sel ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m1_nxt_st[48:0] = S_S0_WAIT;
                  end
       endcase
  end
  S_S1_WAIT:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       case(1'b1)
         ~m1_s1_hld: begin
                          m1_nxt_st[48:0] = m1_s1_wt_sel ? S_S1_GNT : s1_hready ? S_S1_DATA : S_S1_CMD;
                          m1_s1_cmd_last = m1_s1_wt_sel ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m1_nxt_st[48:0] = S_S1_WAIT;
                  end
       endcase
  end
  S_S2_WAIT:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       case(1'b1)
         ~m1_s2_hld: begin
                          m1_nxt_st[48:0] = m1_s2_wt_sel ? S_S2_GNT : s2_hready ? S_S2_DATA : S_S2_CMD;
                          m1_s2_cmd_last = m1_s2_wt_sel ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m1_nxt_st[48:0] = S_S2_WAIT;
                  end
       endcase
  end
  S_S3_WAIT:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       case(1'b1)
         ~m1_s3_hld: begin
                          m1_nxt_st[48:0] = m1_s3_wt_sel ? S_S3_GNT : s3_hready ? S_S3_DATA : S_S3_CMD;
                          m1_s3_cmd_last = m1_s3_wt_sel ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m1_nxt_st[48:0] = S_S3_WAIT;
                  end
       endcase
  end
  S_S4_WAIT:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       case(1'b1)
         ~m1_s4_hld: begin
                          m1_nxt_st[48:0] = m1_s4_wt_sel ? S_S4_GNT : s4_hready ? S_S4_DATA : S_S4_CMD;
                          m1_s4_cmd_last = m1_s4_wt_sel ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m1_nxt_st[48:0] = S_S4_WAIT;
                  end
       endcase
  end
  S_S5_WAIT:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       case(1'b1)
         ~m1_s5_hld: begin
                          m1_nxt_st[48:0] = m1_s5_wt_sel ? S_S5_GNT : s5_hready ? S_S5_DATA : S_S5_CMD;
                          m1_s5_cmd_last = m1_s5_wt_sel ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m1_nxt_st[48:0] = S_S5_WAIT;
                  end
       endcase
  end
  S_S6_WAIT:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       case(1'b1)
         ~m1_s6_hld: begin
                          m1_nxt_st[48:0] = m1_s6_wt_sel ? S_S6_GNT : s6_hready ? S_S6_DATA : S_S6_CMD;
                          m1_s6_cmd_last = m1_s6_wt_sel ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m1_nxt_st[48:0] = S_S6_WAIT;
                  end
       endcase
  end
  S_S7_WAIT:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       case(1'b1)
         ~m1_s7_hld: begin
                          m1_nxt_st[48:0] = m1_s7_wt_sel ? S_S7_GNT : s7_hready ? S_S7_DATA : S_S7_CMD;
                          m1_s7_cmd_last = m1_s7_wt_sel ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m1_nxt_st[48:0] = S_S7_WAIT;
                  end
       endcase
  end
  S_S8_WAIT:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       case(1'b1)
         ~m1_s8_hld: begin
                          m1_nxt_st[48:0] = m1_s8_wt_sel ? S_S8_GNT : s8_hready ? S_S8_DATA : S_S8_CMD;
                          m1_s8_cmd_last = m1_s8_wt_sel ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m1_nxt_st[48:0] = S_S8_WAIT;
                  end
       endcase
  end
  S_S9_WAIT:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       case(1'b1)
         ~m1_s9_hld: begin
                          m1_nxt_st[48:0] = m1_s9_wt_sel ? S_S9_GNT : s9_hready ? S_S9_DATA : S_S9_CMD;
                          m1_s9_cmd_last = m1_s9_wt_sel ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m1_nxt_st[48:0] = S_S9_WAIT;
                  end
       endcase
  end
  S_S10_WAIT:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       case(1'b1)
         ~m1_s10_hld: begin
                          m1_nxt_st[48:0] = m1_s10_wt_sel ? S_S10_GNT : s10_hready ? S_S10_DATA : S_S10_CMD;
                          m1_s10_cmd_last = m1_s10_wt_sel ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m1_nxt_st[48:0] = S_S10_WAIT;
                  end
       endcase
  end
  S_S11_WAIT:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       case(1'b1)
         ~m1_s11_hld: begin
                          m1_nxt_st[48:0] = m1_s11_wt_sel ? S_S11_GNT : s11_hready ? S_S11_DATA : S_S11_CMD;
                          m1_s11_cmd_last = m1_s11_wt_sel ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m1_nxt_st[48:0] = S_S11_WAIT;
                  end
       endcase
  end
  S_S0_CMD: begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = s0_hready ? 1'b1 : 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       m1_nxt_st[48:0] = s0_hready  ? S_S0_DATA : S_S0_CMD;
  end
  S_S0_DATA:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b1;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       if(s0_hready)
         begin
           case(1'b1)
             m1_s0_sel: begin
                              m1_nxt_st[48:0] = S_S0_DATA;
                              m1_s0_cmd_cur = 1'b1;
                             end
             m1_s0_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S0_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s1_sel: begin
                              m1_nxt_st[48:0] = m1_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m1_latch_cmd = m1_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m1_s1_cmd_cur = m1_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m1_s1_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S1_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s2_sel: begin
                              m1_nxt_st[48:0] = m1_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m1_latch_cmd = m1_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m1_s2_cmd_cur = m1_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m1_s2_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S2_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s3_sel: begin
                              m1_nxt_st[48:0] = m1_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m1_latch_cmd = m1_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m1_s3_cmd_cur = m1_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m1_s3_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S3_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s4_sel: begin
                              m1_nxt_st[48:0] = m1_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m1_latch_cmd = m1_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m1_s4_cmd_cur = m1_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m1_s4_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S4_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s5_sel: begin
                              m1_nxt_st[48:0] = m1_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m1_latch_cmd = m1_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m1_s5_cmd_cur = m1_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m1_s5_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S5_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s6_sel: begin
                              m1_nxt_st[48:0] = m1_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m1_latch_cmd = m1_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m1_s6_cmd_cur = m1_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m1_s6_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S6_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s7_sel: begin
                              m1_nxt_st[48:0] = m1_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m1_latch_cmd = m1_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m1_s7_cmd_cur = m1_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m1_s7_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S7_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s8_sel: begin
                              m1_nxt_st[48:0] = m1_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m1_latch_cmd = m1_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m1_s8_cmd_cur = m1_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m1_s8_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S8_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s9_sel: begin
                              m1_nxt_st[48:0] = m1_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m1_latch_cmd = m1_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m1_s9_cmd_cur = m1_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m1_s9_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S9_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s10_sel: begin
                              m1_nxt_st[48:0] = m1_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m1_latch_cmd = m1_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m1_s10_cmd_cur = m1_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m1_s10_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S10_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s11_sel: begin
                              m1_nxt_st[48:0] = m1_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m1_latch_cmd = m1_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m1_s11_cmd_cur = m1_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m1_s11_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S11_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             default: begin
                             m1_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m1_nxt_st[48:0] = S_S0_DATA;
end
  S_S1_CMD: begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = s1_hready ? 1'b1 : 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       m1_nxt_st[48:0] = s1_hready  ? S_S1_DATA : S_S1_CMD;
  end
  S_S1_DATA:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b1;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       if(s1_hready)
         begin
           case(1'b1)
             m1_s0_sel: begin
                              m1_nxt_st[48:0] = m1_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m1_latch_cmd = m1_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m1_s0_cmd_cur = m1_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m1_s0_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S0_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s1_sel: begin
                              m1_nxt_st[48:0] = S_S1_DATA;
                              m1_s1_cmd_cur = 1'b1;
                             end
             m1_s1_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S1_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s2_sel: begin
                              m1_nxt_st[48:0] = m1_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m1_latch_cmd = m1_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m1_s2_cmd_cur = m1_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m1_s2_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S2_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s3_sel: begin
                              m1_nxt_st[48:0] = m1_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m1_latch_cmd = m1_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m1_s3_cmd_cur = m1_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m1_s3_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S3_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s4_sel: begin
                              m1_nxt_st[48:0] = m1_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m1_latch_cmd = m1_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m1_s4_cmd_cur = m1_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m1_s4_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S4_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s5_sel: begin
                              m1_nxt_st[48:0] = m1_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m1_latch_cmd = m1_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m1_s5_cmd_cur = m1_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m1_s5_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S5_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s6_sel: begin
                              m1_nxt_st[48:0] = m1_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m1_latch_cmd = m1_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m1_s6_cmd_cur = m1_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m1_s6_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S6_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s7_sel: begin
                              m1_nxt_st[48:0] = m1_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m1_latch_cmd = m1_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m1_s7_cmd_cur = m1_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m1_s7_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S7_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s8_sel: begin
                              m1_nxt_st[48:0] = m1_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m1_latch_cmd = m1_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m1_s8_cmd_cur = m1_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m1_s8_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S8_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s9_sel: begin
                              m1_nxt_st[48:0] = m1_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m1_latch_cmd = m1_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m1_s9_cmd_cur = m1_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m1_s9_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S9_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s10_sel: begin
                              m1_nxt_st[48:0] = m1_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m1_latch_cmd = m1_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m1_s10_cmd_cur = m1_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m1_s10_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S10_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s11_sel: begin
                              m1_nxt_st[48:0] = m1_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m1_latch_cmd = m1_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m1_s11_cmd_cur = m1_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m1_s11_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S11_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             default: begin
                             m1_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m1_nxt_st[48:0] = S_S1_DATA;
end
  S_S2_CMD: begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = s2_hready ? 1'b1 : 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       m1_nxt_st[48:0] = s2_hready  ? S_S2_DATA : S_S2_CMD;
  end
  S_S2_DATA:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b1;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       if(s2_hready)
         begin
           case(1'b1)
             m1_s0_sel: begin
                              m1_nxt_st[48:0] = m1_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m1_latch_cmd = m1_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m1_s0_cmd_cur = m1_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m1_s0_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S0_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s1_sel: begin
                              m1_nxt_st[48:0] = m1_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m1_latch_cmd = m1_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m1_s1_cmd_cur = m1_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m1_s1_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S1_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s2_sel: begin
                              m1_nxt_st[48:0] = S_S2_DATA;
                              m1_s2_cmd_cur = 1'b1;
                             end
             m1_s2_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S2_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s3_sel: begin
                              m1_nxt_st[48:0] = m1_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m1_latch_cmd = m1_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m1_s3_cmd_cur = m1_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m1_s3_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S3_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s4_sel: begin
                              m1_nxt_st[48:0] = m1_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m1_latch_cmd = m1_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m1_s4_cmd_cur = m1_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m1_s4_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S4_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s5_sel: begin
                              m1_nxt_st[48:0] = m1_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m1_latch_cmd = m1_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m1_s5_cmd_cur = m1_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m1_s5_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S5_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s6_sel: begin
                              m1_nxt_st[48:0] = m1_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m1_latch_cmd = m1_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m1_s6_cmd_cur = m1_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m1_s6_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S6_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s7_sel: begin
                              m1_nxt_st[48:0] = m1_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m1_latch_cmd = m1_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m1_s7_cmd_cur = m1_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m1_s7_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S7_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s8_sel: begin
                              m1_nxt_st[48:0] = m1_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m1_latch_cmd = m1_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m1_s8_cmd_cur = m1_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m1_s8_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S8_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s9_sel: begin
                              m1_nxt_st[48:0] = m1_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m1_latch_cmd = m1_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m1_s9_cmd_cur = m1_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m1_s9_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S9_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s10_sel: begin
                              m1_nxt_st[48:0] = m1_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m1_latch_cmd = m1_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m1_s10_cmd_cur = m1_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m1_s10_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S10_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s11_sel: begin
                              m1_nxt_st[48:0] = m1_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m1_latch_cmd = m1_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m1_s11_cmd_cur = m1_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m1_s11_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S11_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             default: begin
                             m1_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m1_nxt_st[48:0] = S_S2_DATA;
end
  S_S3_CMD: begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = s3_hready ? 1'b1 : 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       m1_nxt_st[48:0] = s3_hready  ? S_S3_DATA : S_S3_CMD;
  end
  S_S3_DATA:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b1;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       if(s3_hready)
         begin
           case(1'b1)
             m1_s0_sel: begin
                              m1_nxt_st[48:0] = m1_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m1_latch_cmd = m1_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m1_s0_cmd_cur = m1_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m1_s0_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S0_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s1_sel: begin
                              m1_nxt_st[48:0] = m1_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m1_latch_cmd = m1_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m1_s1_cmd_cur = m1_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m1_s1_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S1_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s2_sel: begin
                              m1_nxt_st[48:0] = m1_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m1_latch_cmd = m1_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m1_s2_cmd_cur = m1_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m1_s2_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S2_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s3_sel: begin
                              m1_nxt_st[48:0] = S_S3_DATA;
                              m1_s3_cmd_cur = 1'b1;
                             end
             m1_s3_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S3_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s4_sel: begin
                              m1_nxt_st[48:0] = m1_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m1_latch_cmd = m1_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m1_s4_cmd_cur = m1_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m1_s4_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S4_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s5_sel: begin
                              m1_nxt_st[48:0] = m1_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m1_latch_cmd = m1_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m1_s5_cmd_cur = m1_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m1_s5_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S5_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s6_sel: begin
                              m1_nxt_st[48:0] = m1_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m1_latch_cmd = m1_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m1_s6_cmd_cur = m1_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m1_s6_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S6_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s7_sel: begin
                              m1_nxt_st[48:0] = m1_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m1_latch_cmd = m1_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m1_s7_cmd_cur = m1_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m1_s7_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S7_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s8_sel: begin
                              m1_nxt_st[48:0] = m1_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m1_latch_cmd = m1_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m1_s8_cmd_cur = m1_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m1_s8_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S8_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s9_sel: begin
                              m1_nxt_st[48:0] = m1_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m1_latch_cmd = m1_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m1_s9_cmd_cur = m1_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m1_s9_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S9_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s10_sel: begin
                              m1_nxt_st[48:0] = m1_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m1_latch_cmd = m1_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m1_s10_cmd_cur = m1_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m1_s10_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S10_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s11_sel: begin
                              m1_nxt_st[48:0] = m1_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m1_latch_cmd = m1_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m1_s11_cmd_cur = m1_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m1_s11_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S11_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             default: begin
                             m1_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m1_nxt_st[48:0] = S_S3_DATA;
end
  S_S4_CMD: begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = s4_hready ? 1'b1 : 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       m1_nxt_st[48:0] = s4_hready  ? S_S4_DATA : S_S4_CMD;
  end
  S_S4_DATA:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b1;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       if(s4_hready)
         begin
           case(1'b1)
             m1_s0_sel: begin
                              m1_nxt_st[48:0] = m1_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m1_latch_cmd = m1_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m1_s0_cmd_cur = m1_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m1_s0_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S0_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s1_sel: begin
                              m1_nxt_st[48:0] = m1_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m1_latch_cmd = m1_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m1_s1_cmd_cur = m1_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m1_s1_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S1_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s2_sel: begin
                              m1_nxt_st[48:0] = m1_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m1_latch_cmd = m1_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m1_s2_cmd_cur = m1_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m1_s2_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S2_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s3_sel: begin
                              m1_nxt_st[48:0] = m1_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m1_latch_cmd = m1_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m1_s3_cmd_cur = m1_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m1_s3_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S3_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s4_sel: begin
                              m1_nxt_st[48:0] = S_S4_DATA;
                              m1_s4_cmd_cur = 1'b1;
                             end
             m1_s4_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S4_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s5_sel: begin
                              m1_nxt_st[48:0] = m1_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m1_latch_cmd = m1_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m1_s5_cmd_cur = m1_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m1_s5_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S5_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s6_sel: begin
                              m1_nxt_st[48:0] = m1_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m1_latch_cmd = m1_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m1_s6_cmd_cur = m1_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m1_s6_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S6_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s7_sel: begin
                              m1_nxt_st[48:0] = m1_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m1_latch_cmd = m1_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m1_s7_cmd_cur = m1_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m1_s7_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S7_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s8_sel: begin
                              m1_nxt_st[48:0] = m1_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m1_latch_cmd = m1_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m1_s8_cmd_cur = m1_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m1_s8_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S8_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s9_sel: begin
                              m1_nxt_st[48:0] = m1_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m1_latch_cmd = m1_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m1_s9_cmd_cur = m1_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m1_s9_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S9_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s10_sel: begin
                              m1_nxt_st[48:0] = m1_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m1_latch_cmd = m1_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m1_s10_cmd_cur = m1_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m1_s10_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S10_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s11_sel: begin
                              m1_nxt_st[48:0] = m1_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m1_latch_cmd = m1_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m1_s11_cmd_cur = m1_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m1_s11_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S11_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             default: begin
                             m1_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m1_nxt_st[48:0] = S_S4_DATA;
end
  S_S5_CMD: begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = s5_hready ? 1'b1 : 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       m1_nxt_st[48:0] = s5_hready  ? S_S5_DATA : S_S5_CMD;
  end
  S_S5_DATA:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b1;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       if(s5_hready)
         begin
           case(1'b1)
             m1_s0_sel: begin
                              m1_nxt_st[48:0] = m1_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m1_latch_cmd = m1_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m1_s0_cmd_cur = m1_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m1_s0_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S0_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s1_sel: begin
                              m1_nxt_st[48:0] = m1_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m1_latch_cmd = m1_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m1_s1_cmd_cur = m1_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m1_s1_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S1_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s2_sel: begin
                              m1_nxt_st[48:0] = m1_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m1_latch_cmd = m1_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m1_s2_cmd_cur = m1_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m1_s2_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S2_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s3_sel: begin
                              m1_nxt_st[48:0] = m1_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m1_latch_cmd = m1_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m1_s3_cmd_cur = m1_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m1_s3_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S3_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s4_sel: begin
                              m1_nxt_st[48:0] = m1_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m1_latch_cmd = m1_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m1_s4_cmd_cur = m1_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m1_s4_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S4_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s5_sel: begin
                              m1_nxt_st[48:0] = S_S5_DATA;
                              m1_s5_cmd_cur = 1'b1;
                             end
             m1_s5_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S5_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s6_sel: begin
                              m1_nxt_st[48:0] = m1_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m1_latch_cmd = m1_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m1_s6_cmd_cur = m1_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m1_s6_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S6_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s7_sel: begin
                              m1_nxt_st[48:0] = m1_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m1_latch_cmd = m1_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m1_s7_cmd_cur = m1_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m1_s7_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S7_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s8_sel: begin
                              m1_nxt_st[48:0] = m1_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m1_latch_cmd = m1_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m1_s8_cmd_cur = m1_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m1_s8_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S8_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s9_sel: begin
                              m1_nxt_st[48:0] = m1_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m1_latch_cmd = m1_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m1_s9_cmd_cur = m1_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m1_s9_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S9_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s10_sel: begin
                              m1_nxt_st[48:0] = m1_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m1_latch_cmd = m1_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m1_s10_cmd_cur = m1_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m1_s10_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S10_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s11_sel: begin
                              m1_nxt_st[48:0] = m1_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m1_latch_cmd = m1_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m1_s11_cmd_cur = m1_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m1_s11_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S11_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             default: begin
                             m1_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m1_nxt_st[48:0] = S_S5_DATA;
end
  S_S6_CMD: begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = s6_hready ? 1'b1 : 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       m1_nxt_st[48:0] = s6_hready  ? S_S6_DATA : S_S6_CMD;
  end
  S_S6_DATA:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b1;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       if(s6_hready)
         begin
           case(1'b1)
             m1_s0_sel: begin
                              m1_nxt_st[48:0] = m1_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m1_latch_cmd = m1_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m1_s0_cmd_cur = m1_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m1_s0_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S0_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s1_sel: begin
                              m1_nxt_st[48:0] = m1_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m1_latch_cmd = m1_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m1_s1_cmd_cur = m1_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m1_s1_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S1_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s2_sel: begin
                              m1_nxt_st[48:0] = m1_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m1_latch_cmd = m1_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m1_s2_cmd_cur = m1_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m1_s2_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S2_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s3_sel: begin
                              m1_nxt_st[48:0] = m1_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m1_latch_cmd = m1_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m1_s3_cmd_cur = m1_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m1_s3_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S3_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s4_sel: begin
                              m1_nxt_st[48:0] = m1_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m1_latch_cmd = m1_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m1_s4_cmd_cur = m1_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m1_s4_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S4_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s5_sel: begin
                              m1_nxt_st[48:0] = m1_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m1_latch_cmd = m1_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m1_s5_cmd_cur = m1_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m1_s5_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S5_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s6_sel: begin
                              m1_nxt_st[48:0] = S_S6_DATA;
                              m1_s6_cmd_cur = 1'b1;
                             end
             m1_s6_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S6_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s7_sel: begin
                              m1_nxt_st[48:0] = m1_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m1_latch_cmd = m1_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m1_s7_cmd_cur = m1_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m1_s7_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S7_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s8_sel: begin
                              m1_nxt_st[48:0] = m1_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m1_latch_cmd = m1_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m1_s8_cmd_cur = m1_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m1_s8_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S8_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s9_sel: begin
                              m1_nxt_st[48:0] = m1_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m1_latch_cmd = m1_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m1_s9_cmd_cur = m1_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m1_s9_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S9_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s10_sel: begin
                              m1_nxt_st[48:0] = m1_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m1_latch_cmd = m1_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m1_s10_cmd_cur = m1_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m1_s10_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S10_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s11_sel: begin
                              m1_nxt_st[48:0] = m1_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m1_latch_cmd = m1_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m1_s11_cmd_cur = m1_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m1_s11_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S11_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             default: begin
                             m1_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m1_nxt_st[48:0] = S_S6_DATA;
end
  S_S7_CMD: begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = s7_hready ? 1'b1 : 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       m1_nxt_st[48:0] = s7_hready  ? S_S7_DATA : S_S7_CMD;
  end
  S_S7_DATA:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b1;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       if(s7_hready)
         begin
           case(1'b1)
             m1_s0_sel: begin
                              m1_nxt_st[48:0] = m1_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m1_latch_cmd = m1_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m1_s0_cmd_cur = m1_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m1_s0_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S0_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s1_sel: begin
                              m1_nxt_st[48:0] = m1_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m1_latch_cmd = m1_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m1_s1_cmd_cur = m1_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m1_s1_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S1_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s2_sel: begin
                              m1_nxt_st[48:0] = m1_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m1_latch_cmd = m1_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m1_s2_cmd_cur = m1_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m1_s2_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S2_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s3_sel: begin
                              m1_nxt_st[48:0] = m1_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m1_latch_cmd = m1_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m1_s3_cmd_cur = m1_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m1_s3_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S3_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s4_sel: begin
                              m1_nxt_st[48:0] = m1_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m1_latch_cmd = m1_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m1_s4_cmd_cur = m1_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m1_s4_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S4_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s5_sel: begin
                              m1_nxt_st[48:0] = m1_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m1_latch_cmd = m1_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m1_s5_cmd_cur = m1_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m1_s5_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S5_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s6_sel: begin
                              m1_nxt_st[48:0] = m1_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m1_latch_cmd = m1_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m1_s6_cmd_cur = m1_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m1_s6_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S6_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s7_sel: begin
                              m1_nxt_st[48:0] = S_S7_DATA;
                              m1_s7_cmd_cur = 1'b1;
                             end
             m1_s7_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S7_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s8_sel: begin
                              m1_nxt_st[48:0] = m1_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m1_latch_cmd = m1_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m1_s8_cmd_cur = m1_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m1_s8_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S8_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s9_sel: begin
                              m1_nxt_st[48:0] = m1_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m1_latch_cmd = m1_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m1_s9_cmd_cur = m1_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m1_s9_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S9_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s10_sel: begin
                              m1_nxt_st[48:0] = m1_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m1_latch_cmd = m1_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m1_s10_cmd_cur = m1_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m1_s10_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S10_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s11_sel: begin
                              m1_nxt_st[48:0] = m1_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m1_latch_cmd = m1_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m1_s11_cmd_cur = m1_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m1_s11_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S11_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             default: begin
                             m1_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m1_nxt_st[48:0] = S_S7_DATA;
end
  S_S8_CMD: begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = s8_hready ? 1'b1 : 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       m1_nxt_st[48:0] = s8_hready  ? S_S8_DATA : S_S8_CMD;
  end
  S_S8_DATA:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b1;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       if(s8_hready)
         begin
           case(1'b1)
             m1_s0_sel: begin
                              m1_nxt_st[48:0] = m1_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m1_latch_cmd = m1_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m1_s0_cmd_cur = m1_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m1_s0_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S0_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s1_sel: begin
                              m1_nxt_st[48:0] = m1_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m1_latch_cmd = m1_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m1_s1_cmd_cur = m1_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m1_s1_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S1_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s2_sel: begin
                              m1_nxt_st[48:0] = m1_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m1_latch_cmd = m1_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m1_s2_cmd_cur = m1_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m1_s2_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S2_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s3_sel: begin
                              m1_nxt_st[48:0] = m1_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m1_latch_cmd = m1_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m1_s3_cmd_cur = m1_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m1_s3_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S3_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s4_sel: begin
                              m1_nxt_st[48:0] = m1_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m1_latch_cmd = m1_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m1_s4_cmd_cur = m1_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m1_s4_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S4_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s5_sel: begin
                              m1_nxt_st[48:0] = m1_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m1_latch_cmd = m1_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m1_s5_cmd_cur = m1_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m1_s5_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S5_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s6_sel: begin
                              m1_nxt_st[48:0] = m1_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m1_latch_cmd = m1_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m1_s6_cmd_cur = m1_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m1_s6_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S6_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s7_sel: begin
                              m1_nxt_st[48:0] = m1_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m1_latch_cmd = m1_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m1_s7_cmd_cur = m1_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m1_s7_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S7_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s8_sel: begin
                              m1_nxt_st[48:0] = S_S8_DATA;
                              m1_s8_cmd_cur = 1'b1;
                             end
             m1_s8_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S8_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s9_sel: begin
                              m1_nxt_st[48:0] = m1_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m1_latch_cmd = m1_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m1_s9_cmd_cur = m1_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m1_s9_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S9_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s10_sel: begin
                              m1_nxt_st[48:0] = m1_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m1_latch_cmd = m1_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m1_s10_cmd_cur = m1_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m1_s10_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S10_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s11_sel: begin
                              m1_nxt_st[48:0] = m1_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m1_latch_cmd = m1_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m1_s11_cmd_cur = m1_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m1_s11_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S11_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             default: begin
                             m1_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m1_nxt_st[48:0] = S_S8_DATA;
end
  S_S9_CMD: begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = s9_hready ? 1'b1 : 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       m1_nxt_st[48:0] = s9_hready  ? S_S9_DATA : S_S9_CMD;
  end
  S_S9_DATA:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b1;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       if(s9_hready)
         begin
           case(1'b1)
             m1_s0_sel: begin
                              m1_nxt_st[48:0] = m1_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m1_latch_cmd = m1_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m1_s0_cmd_cur = m1_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m1_s0_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S0_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s1_sel: begin
                              m1_nxt_st[48:0] = m1_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m1_latch_cmd = m1_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m1_s1_cmd_cur = m1_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m1_s1_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S1_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s2_sel: begin
                              m1_nxt_st[48:0] = m1_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m1_latch_cmd = m1_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m1_s2_cmd_cur = m1_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m1_s2_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S2_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s3_sel: begin
                              m1_nxt_st[48:0] = m1_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m1_latch_cmd = m1_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m1_s3_cmd_cur = m1_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m1_s3_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S3_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s4_sel: begin
                              m1_nxt_st[48:0] = m1_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m1_latch_cmd = m1_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m1_s4_cmd_cur = m1_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m1_s4_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S4_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s5_sel: begin
                              m1_nxt_st[48:0] = m1_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m1_latch_cmd = m1_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m1_s5_cmd_cur = m1_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m1_s5_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S5_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s6_sel: begin
                              m1_nxt_st[48:0] = m1_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m1_latch_cmd = m1_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m1_s6_cmd_cur = m1_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m1_s6_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S6_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s7_sel: begin
                              m1_nxt_st[48:0] = m1_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m1_latch_cmd = m1_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m1_s7_cmd_cur = m1_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m1_s7_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S7_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s8_sel: begin
                              m1_nxt_st[48:0] = m1_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m1_latch_cmd = m1_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m1_s8_cmd_cur = m1_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m1_s8_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S8_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s9_sel: begin
                              m1_nxt_st[48:0] = S_S9_DATA;
                              m1_s9_cmd_cur = 1'b1;
                             end
             m1_s9_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S9_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s10_sel: begin
                              m1_nxt_st[48:0] = m1_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m1_latch_cmd = m1_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m1_s10_cmd_cur = m1_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m1_s10_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S10_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s11_sel: begin
                              m1_nxt_st[48:0] = m1_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m1_latch_cmd = m1_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m1_s11_cmd_cur = m1_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m1_s11_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S11_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             default: begin
                             m1_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m1_nxt_st[48:0] = S_S9_DATA;
end
  S_S10_CMD: begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = s10_hready ? 1'b1 : 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       m1_nxt_st[48:0] = s10_hready  ? S_S10_DATA : S_S10_CMD;
  end
  S_S10_DATA:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b1;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       if(s10_hready)
         begin
           case(1'b1)
             m1_s0_sel: begin
                              m1_nxt_st[48:0] = m1_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m1_latch_cmd = m1_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m1_s0_cmd_cur = m1_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m1_s0_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S0_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s1_sel: begin
                              m1_nxt_st[48:0] = m1_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m1_latch_cmd = m1_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m1_s1_cmd_cur = m1_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m1_s1_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S1_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s2_sel: begin
                              m1_nxt_st[48:0] = m1_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m1_latch_cmd = m1_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m1_s2_cmd_cur = m1_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m1_s2_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S2_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s3_sel: begin
                              m1_nxt_st[48:0] = m1_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m1_latch_cmd = m1_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m1_s3_cmd_cur = m1_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m1_s3_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S3_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s4_sel: begin
                              m1_nxt_st[48:0] = m1_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m1_latch_cmd = m1_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m1_s4_cmd_cur = m1_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m1_s4_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S4_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s5_sel: begin
                              m1_nxt_st[48:0] = m1_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m1_latch_cmd = m1_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m1_s5_cmd_cur = m1_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m1_s5_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S5_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s6_sel: begin
                              m1_nxt_st[48:0] = m1_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m1_latch_cmd = m1_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m1_s6_cmd_cur = m1_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m1_s6_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S6_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s7_sel: begin
                              m1_nxt_st[48:0] = m1_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m1_latch_cmd = m1_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m1_s7_cmd_cur = m1_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m1_s7_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S7_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s8_sel: begin
                              m1_nxt_st[48:0] = m1_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m1_latch_cmd = m1_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m1_s8_cmd_cur = m1_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m1_s8_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S8_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s9_sel: begin
                              m1_nxt_st[48:0] = m1_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m1_latch_cmd = m1_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m1_s9_cmd_cur = m1_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m1_s9_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S9_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s10_sel: begin
                              m1_nxt_st[48:0] = S_S10_DATA;
                              m1_s10_cmd_cur = 1'b1;
                             end
             m1_s10_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S10_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s11_sel: begin
                              m1_nxt_st[48:0] = m1_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m1_latch_cmd = m1_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m1_s11_cmd_cur = m1_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m1_s11_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S11_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             default: begin
                             m1_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m1_nxt_st[48:0] = S_S10_DATA;
end
  S_S11_CMD: begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = s11_hready ? 1'b1 : 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b0;
       m1_nxt_st[48:0] = s11_hready  ? S_S11_DATA : S_S11_CMD;
  end
  S_S11_DATA:begin
       m1_latch_cmd = 1'b0;
       m1_s0_cmd_last = 1'b0;
       m1_s0_cmd_cur = 1'b0;
       m1_s0_data = 1'b0;
       m1_s1_cmd_last = 1'b0;
       m1_s1_cmd_cur = 1'b0;
       m1_s1_data = 1'b0;
       m1_s2_cmd_last = 1'b0;
       m1_s2_cmd_cur = 1'b0;
       m1_s2_data = 1'b0;
       m1_s3_cmd_last = 1'b0;
       m1_s3_cmd_cur = 1'b0;
       m1_s3_data = 1'b0;
       m1_s4_cmd_last = 1'b0;
       m1_s4_cmd_cur = 1'b0;
       m1_s4_data = 1'b0;
       m1_s5_cmd_last = 1'b0;
       m1_s5_cmd_cur = 1'b0;
       m1_s5_data = 1'b0;
       m1_s6_cmd_last = 1'b0;
       m1_s6_cmd_cur = 1'b0;
       m1_s6_data = 1'b0;
       m1_s7_cmd_last = 1'b0;
       m1_s7_cmd_cur = 1'b0;
       m1_s7_data = 1'b0;
       m1_s8_cmd_last = 1'b0;
       m1_s8_cmd_cur = 1'b0;
       m1_s8_data = 1'b0;
       m1_s9_cmd_last = 1'b0;
       m1_s9_cmd_cur = 1'b0;
       m1_s9_data = 1'b0;
       m1_s10_cmd_last = 1'b0;
       m1_s10_cmd_cur = 1'b0;
       m1_s10_data = 1'b0;
       m1_s11_cmd_last = 1'b0;
       m1_s11_cmd_cur = 1'b0;
       m1_s11_data = 1'b1;
       if(s11_hready)
         begin
           case(1'b1)
             m1_s0_sel: begin
                              m1_nxt_st[48:0] = m1_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m1_latch_cmd = m1_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m1_s0_cmd_cur = m1_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m1_s0_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S0_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s1_sel: begin
                              m1_nxt_st[48:0] = m1_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m1_latch_cmd = m1_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m1_s1_cmd_cur = m1_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m1_s1_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S1_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s2_sel: begin
                              m1_nxt_st[48:0] = m1_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m1_latch_cmd = m1_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m1_s2_cmd_cur = m1_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m1_s2_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S2_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s3_sel: begin
                              m1_nxt_st[48:0] = m1_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m1_latch_cmd = m1_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m1_s3_cmd_cur = m1_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m1_s3_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S3_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s4_sel: begin
                              m1_nxt_st[48:0] = m1_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m1_latch_cmd = m1_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m1_s4_cmd_cur = m1_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m1_s4_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S4_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s5_sel: begin
                              m1_nxt_st[48:0] = m1_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m1_latch_cmd = m1_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m1_s5_cmd_cur = m1_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m1_s5_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S5_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s6_sel: begin
                              m1_nxt_st[48:0] = m1_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m1_latch_cmd = m1_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m1_s6_cmd_cur = m1_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m1_s6_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S6_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s7_sel: begin
                              m1_nxt_st[48:0] = m1_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m1_latch_cmd = m1_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m1_s7_cmd_cur = m1_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m1_s7_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S7_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s8_sel: begin
                              m1_nxt_st[48:0] = m1_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m1_latch_cmd = m1_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m1_s8_cmd_cur = m1_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m1_s8_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S8_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s9_sel: begin
                              m1_nxt_st[48:0] = m1_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m1_latch_cmd = m1_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m1_s9_cmd_cur = m1_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m1_s9_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S9_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s10_sel: begin
                              m1_nxt_st[48:0] = m1_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m1_latch_cmd = m1_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m1_s10_cmd_cur = m1_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m1_s10_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S10_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             m1_s11_sel: begin
                              m1_nxt_st[48:0] = S_S11_DATA;
                              m1_s11_cmd_cur = 1'b1;
                             end
             m1_s11_wt_sel: begin
                                 m1_nxt_st[48:0] = S_S11_GNT;
                                 m1_latch_cmd = 1'b1;
                               end
             default: begin
                             m1_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m1_nxt_st[48:0] = S_S11_DATA;
end
  default: begin
             m1_latch_cmd = 1'b0;
             m1_s0_cmd_last = 1'b0;
             m1_s0_cmd_cur = 1'b0;
             m1_s0_data = 1'b0;
             m1_s1_cmd_last = 1'b0;
             m1_s1_cmd_cur = 1'b0;
             m1_s1_data = 1'b0;
             m1_s2_cmd_last = 1'b0;
             m1_s2_cmd_cur = 1'b0;
             m1_s2_data = 1'b0;
             m1_s3_cmd_last = 1'b0;
             m1_s3_cmd_cur = 1'b0;
             m1_s3_data = 1'b0;
             m1_s4_cmd_last = 1'b0;
             m1_s4_cmd_cur = 1'b0;
             m1_s4_data = 1'b0;
             m1_s5_cmd_last = 1'b0;
             m1_s5_cmd_cur = 1'b0;
             m1_s5_data = 1'b0;
             m1_s6_cmd_last = 1'b0;
             m1_s6_cmd_cur = 1'b0;
             m1_s6_data = 1'b0;
             m1_s7_cmd_last = 1'b0;
             m1_s7_cmd_cur = 1'b0;
             m1_s7_data = 1'b0;
             m1_s8_cmd_last = 1'b0;
             m1_s8_cmd_cur = 1'b0;
             m1_s8_data = 1'b0;
             m1_s9_cmd_last = 1'b0;
             m1_s9_cmd_cur = 1'b0;
             m1_s9_data = 1'b0;
             m1_s10_cmd_last = 1'b0;
             m1_s10_cmd_cur = 1'b0;
             m1_s10_data = 1'b0;
             m1_s11_cmd_last = 1'b0;
             m1_s11_cmd_cur = 1'b0;
             m1_s11_data = 1'b0;
             m1_nxt_st[48:0] = S_IDLE;
  end
endcase
end
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
       m2_cur_st[48:0] <= S_IDLE;
    else
       m2_cur_st[48:0] <= m2_nxt_st[48:0];
  end
always @ (*)
begin
case(m2_cur_st[48:0])
  S_IDLE:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       case(1'b1)
         m2_s0_sel: begin
                          m2_nxt_st[48:0] = m2_s0_hld ? S_S0_WAIT : (s0_hready ? S_S0_DATA : S_S0_CMD);
                          m2_latch_cmd = m2_s0_hld ? 1'b1 : (s0_hready ? 1'b0 : 1'b1);
                          m2_s0_cmd_cur = m2_s0_hld ? 1'b0 : (s0_hready ? 1'b1 : 1'b0);
                        end
         m2_s0_wt_sel: begin
                             m2_nxt_st[48:0] = S_S0_GNT;
                             m2_latch_cmd = 1'b1;
                           end
         m2_s1_sel: begin
                          m2_nxt_st[48:0] = m2_s1_hld ? S_S1_WAIT : (s1_hready ? S_S1_DATA : S_S1_CMD);
                          m2_latch_cmd = m2_s1_hld ? 1'b1 : (s1_hready ? 1'b0 : 1'b1);
                          m2_s1_cmd_cur = m2_s1_hld ? 1'b0 : (s1_hready ? 1'b1 : 1'b0);
                        end
         m2_s1_wt_sel: begin
                             m2_nxt_st[48:0] = S_S1_GNT;
                             m2_latch_cmd = 1'b1;
                           end
         m2_s2_sel: begin
                          m2_nxt_st[48:0] = m2_s2_hld ? S_S2_WAIT : (s2_hready ? S_S2_DATA : S_S2_CMD);
                          m2_latch_cmd = m2_s2_hld ? 1'b1 : (s2_hready ? 1'b0 : 1'b1);
                          m2_s2_cmd_cur = m2_s2_hld ? 1'b0 : (s2_hready ? 1'b1 : 1'b0);
                        end
         m2_s2_wt_sel: begin
                             m2_nxt_st[48:0] = S_S2_GNT;
                             m2_latch_cmd = 1'b1;
                           end
         m2_s3_sel: begin
                          m2_nxt_st[48:0] = m2_s3_hld ? S_S3_WAIT : (s3_hready ? S_S3_DATA : S_S3_CMD);
                          m2_latch_cmd = m2_s3_hld ? 1'b1 : (s3_hready ? 1'b0 : 1'b1);
                          m2_s3_cmd_cur = m2_s3_hld ? 1'b0 : (s3_hready ? 1'b1 : 1'b0);
                        end
         m2_s3_wt_sel: begin
                             m2_nxt_st[48:0] = S_S3_GNT;
                             m2_latch_cmd = 1'b1;
                           end
         m2_s4_sel: begin
                          m2_nxt_st[48:0] = m2_s4_hld ? S_S4_WAIT : (s4_hready ? S_S4_DATA : S_S4_CMD);
                          m2_latch_cmd = m2_s4_hld ? 1'b1 : (s4_hready ? 1'b0 : 1'b1);
                          m2_s4_cmd_cur = m2_s4_hld ? 1'b0 : (s4_hready ? 1'b1 : 1'b0);
                        end
         m2_s4_wt_sel: begin
                             m2_nxt_st[48:0] = S_S4_GNT;
                             m2_latch_cmd = 1'b1;
                           end
         m2_s5_sel: begin
                          m2_nxt_st[48:0] = m2_s5_hld ? S_S5_WAIT : (s5_hready ? S_S5_DATA : S_S5_CMD);
                          m2_latch_cmd = m2_s5_hld ? 1'b1 : (s5_hready ? 1'b0 : 1'b1);
                          m2_s5_cmd_cur = m2_s5_hld ? 1'b0 : (s5_hready ? 1'b1 : 1'b0);
                        end
         m2_s5_wt_sel: begin
                             m2_nxt_st[48:0] = S_S5_GNT;
                             m2_latch_cmd = 1'b1;
                           end
         m2_s6_sel: begin
                          m2_nxt_st[48:0] = m2_s6_hld ? S_S6_WAIT : (s6_hready ? S_S6_DATA : S_S6_CMD);
                          m2_latch_cmd = m2_s6_hld ? 1'b1 : (s6_hready ? 1'b0 : 1'b1);
                          m2_s6_cmd_cur = m2_s6_hld ? 1'b0 : (s6_hready ? 1'b1 : 1'b0);
                        end
         m2_s6_wt_sel: begin
                             m2_nxt_st[48:0] = S_S6_GNT;
                             m2_latch_cmd = 1'b1;
                           end
         m2_s7_sel: begin
                          m2_nxt_st[48:0] = m2_s7_hld ? S_S7_WAIT : (s7_hready ? S_S7_DATA : S_S7_CMD);
                          m2_latch_cmd = m2_s7_hld ? 1'b1 : (s7_hready ? 1'b0 : 1'b1);
                          m2_s7_cmd_cur = m2_s7_hld ? 1'b0 : (s7_hready ? 1'b1 : 1'b0);
                        end
         m2_s7_wt_sel: begin
                             m2_nxt_st[48:0] = S_S7_GNT;
                             m2_latch_cmd = 1'b1;
                           end
         m2_s8_sel: begin
                          m2_nxt_st[48:0] = m2_s8_hld ? S_S8_WAIT : (s8_hready ? S_S8_DATA : S_S8_CMD);
                          m2_latch_cmd = m2_s8_hld ? 1'b1 : (s8_hready ? 1'b0 : 1'b1);
                          m2_s8_cmd_cur = m2_s8_hld ? 1'b0 : (s8_hready ? 1'b1 : 1'b0);
                        end
         m2_s8_wt_sel: begin
                             m2_nxt_st[48:0] = S_S8_GNT;
                             m2_latch_cmd = 1'b1;
                           end
         m2_s9_sel: begin
                          m2_nxt_st[48:0] = m2_s9_hld ? S_S9_WAIT : (s9_hready ? S_S9_DATA : S_S9_CMD);
                          m2_latch_cmd = m2_s9_hld ? 1'b1 : (s9_hready ? 1'b0 : 1'b1);
                          m2_s9_cmd_cur = m2_s9_hld ? 1'b0 : (s9_hready ? 1'b1 : 1'b0);
                        end
         m2_s9_wt_sel: begin
                             m2_nxt_st[48:0] = S_S9_GNT;
                             m2_latch_cmd = 1'b1;
                           end
         m2_s10_sel: begin
                          m2_nxt_st[48:0] = m2_s10_hld ? S_S10_WAIT : (s10_hready ? S_S10_DATA : S_S10_CMD);
                          m2_latch_cmd = m2_s10_hld ? 1'b1 : (s10_hready ? 1'b0 : 1'b1);
                          m2_s10_cmd_cur = m2_s10_hld ? 1'b0 : (s10_hready ? 1'b1 : 1'b0);
                        end
         m2_s10_wt_sel: begin
                             m2_nxt_st[48:0] = S_S10_GNT;
                             m2_latch_cmd = 1'b1;
                           end
         m2_s11_sel: begin
                          m2_nxt_st[48:0] = m2_s11_hld ? S_S11_WAIT : (s11_hready ? S_S11_DATA : S_S11_CMD);
                          m2_latch_cmd = m2_s11_hld ? 1'b1 : (s11_hready ? 1'b0 : 1'b1);
                          m2_s11_cmd_cur = m2_s11_hld ? 1'b0 : (s11_hready ? 1'b1 : 1'b0);
                        end
         m2_s11_wt_sel: begin
                             m2_nxt_st[48:0] = S_S11_GNT;
                             m2_latch_cmd = 1'b1;
                           end
         default: begin
                          m2_nxt_st[48:0] = S_IDLE;
                  end
       endcase
  end
  S_S0_GNT:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       case(1'b1)
         m2_s0_sel: begin
                          m2_nxt_st[48:0] = m2_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                          m2_s0_cmd_last = m2_s0_hld ? 1'b0 : (s0_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m2_nxt_st[48:0] = S_S0_GNT;
                  end
       endcase
  end
  S_S1_GNT:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       case(1'b1)
         m2_s1_sel: begin
                          m2_nxt_st[48:0] = m2_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                          m2_s1_cmd_last = m2_s1_hld ? 1'b0 : (s1_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m2_nxt_st[48:0] = S_S1_GNT;
                  end
       endcase
  end
  S_S2_GNT:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       case(1'b1)
         m2_s2_sel: begin
                          m2_nxt_st[48:0] = m2_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                          m2_s2_cmd_last = m2_s2_hld ? 1'b0 : (s2_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m2_nxt_st[48:0] = S_S2_GNT;
                  end
       endcase
  end
  S_S3_GNT:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       case(1'b1)
         m2_s3_sel: begin
                          m2_nxt_st[48:0] = m2_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                          m2_s3_cmd_last = m2_s3_hld ? 1'b0 : (s3_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m2_nxt_st[48:0] = S_S3_GNT;
                  end
       endcase
  end
  S_S4_GNT:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       case(1'b1)
         m2_s4_sel: begin
                          m2_nxt_st[48:0] = m2_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                          m2_s4_cmd_last = m2_s4_hld ? 1'b0 : (s4_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m2_nxt_st[48:0] = S_S4_GNT;
                  end
       endcase
  end
  S_S5_GNT:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       case(1'b1)
         m2_s5_sel: begin
                          m2_nxt_st[48:0] = m2_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                          m2_s5_cmd_last = m2_s5_hld ? 1'b0 : (s5_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m2_nxt_st[48:0] = S_S5_GNT;
                  end
       endcase
  end
  S_S6_GNT:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       case(1'b1)
         m2_s6_sel: begin
                          m2_nxt_st[48:0] = m2_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                          m2_s6_cmd_last = m2_s6_hld ? 1'b0 : (s6_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m2_nxt_st[48:0] = S_S6_GNT;
                  end
       endcase
  end
  S_S7_GNT:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       case(1'b1)
         m2_s7_sel: begin
                          m2_nxt_st[48:0] = m2_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                          m2_s7_cmd_last = m2_s7_hld ? 1'b0 : (s7_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m2_nxt_st[48:0] = S_S7_GNT;
                  end
       endcase
  end
  S_S8_GNT:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       case(1'b1)
         m2_s8_sel: begin
                          m2_nxt_st[48:0] = m2_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                          m2_s8_cmd_last = m2_s8_hld ? 1'b0 : (s8_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m2_nxt_st[48:0] = S_S8_GNT;
                  end
       endcase
  end
  S_S9_GNT:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       case(1'b1)
         m2_s9_sel: begin
                          m2_nxt_st[48:0] = m2_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                          m2_s9_cmd_last = m2_s9_hld ? 1'b0 : (s9_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m2_nxt_st[48:0] = S_S9_GNT;
                  end
       endcase
  end
  S_S10_GNT:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       case(1'b1)
         m2_s10_sel: begin
                          m2_nxt_st[48:0] = m2_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                          m2_s10_cmd_last = m2_s10_hld ? 1'b0 : (s10_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m2_nxt_st[48:0] = S_S10_GNT;
                  end
       endcase
  end
  S_S11_GNT:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       case(1'b1)
         m2_s11_sel: begin
                          m2_nxt_st[48:0] = m2_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                          m2_s11_cmd_last = m2_s11_hld ? 1'b0 : (s11_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m2_nxt_st[48:0] = S_S11_GNT;
                  end
       endcase
  end
  S_S0_WAIT:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       case(1'b1)
         ~m2_s0_hld: begin
                          m2_nxt_st[48:0] = m2_s0_wt_sel ? S_S0_GNT : s0_hready ? S_S0_DATA : S_S0_CMD;
                          m2_s0_cmd_last = m2_s0_wt_sel ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m2_nxt_st[48:0] = S_S0_WAIT;
                  end
       endcase
  end
  S_S1_WAIT:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       case(1'b1)
         ~m2_s1_hld: begin
                          m2_nxt_st[48:0] = m2_s1_wt_sel ? S_S1_GNT : s1_hready ? S_S1_DATA : S_S1_CMD;
                          m2_s1_cmd_last = m2_s1_wt_sel ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m2_nxt_st[48:0] = S_S1_WAIT;
                  end
       endcase
  end
  S_S2_WAIT:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       case(1'b1)
         ~m2_s2_hld: begin
                          m2_nxt_st[48:0] = m2_s2_wt_sel ? S_S2_GNT : s2_hready ? S_S2_DATA : S_S2_CMD;
                          m2_s2_cmd_last = m2_s2_wt_sel ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m2_nxt_st[48:0] = S_S2_WAIT;
                  end
       endcase
  end
  S_S3_WAIT:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       case(1'b1)
         ~m2_s3_hld: begin
                          m2_nxt_st[48:0] = m2_s3_wt_sel ? S_S3_GNT : s3_hready ? S_S3_DATA : S_S3_CMD;
                          m2_s3_cmd_last = m2_s3_wt_sel ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m2_nxt_st[48:0] = S_S3_WAIT;
                  end
       endcase
  end
  S_S4_WAIT:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       case(1'b1)
         ~m2_s4_hld: begin
                          m2_nxt_st[48:0] = m2_s4_wt_sel ? S_S4_GNT : s4_hready ? S_S4_DATA : S_S4_CMD;
                          m2_s4_cmd_last = m2_s4_wt_sel ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m2_nxt_st[48:0] = S_S4_WAIT;
                  end
       endcase
  end
  S_S5_WAIT:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       case(1'b1)
         ~m2_s5_hld: begin
                          m2_nxt_st[48:0] = m2_s5_wt_sel ? S_S5_GNT : s5_hready ? S_S5_DATA : S_S5_CMD;
                          m2_s5_cmd_last = m2_s5_wt_sel ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m2_nxt_st[48:0] = S_S5_WAIT;
                  end
       endcase
  end
  S_S6_WAIT:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       case(1'b1)
         ~m2_s6_hld: begin
                          m2_nxt_st[48:0] = m2_s6_wt_sel ? S_S6_GNT : s6_hready ? S_S6_DATA : S_S6_CMD;
                          m2_s6_cmd_last = m2_s6_wt_sel ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m2_nxt_st[48:0] = S_S6_WAIT;
                  end
       endcase
  end
  S_S7_WAIT:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       case(1'b1)
         ~m2_s7_hld: begin
                          m2_nxt_st[48:0] = m2_s7_wt_sel ? S_S7_GNT : s7_hready ? S_S7_DATA : S_S7_CMD;
                          m2_s7_cmd_last = m2_s7_wt_sel ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m2_nxt_st[48:0] = S_S7_WAIT;
                  end
       endcase
  end
  S_S8_WAIT:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       case(1'b1)
         ~m2_s8_hld: begin
                          m2_nxt_st[48:0] = m2_s8_wt_sel ? S_S8_GNT : s8_hready ? S_S8_DATA : S_S8_CMD;
                          m2_s8_cmd_last = m2_s8_wt_sel ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m2_nxt_st[48:0] = S_S8_WAIT;
                  end
       endcase
  end
  S_S9_WAIT:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       case(1'b1)
         ~m2_s9_hld: begin
                          m2_nxt_st[48:0] = m2_s9_wt_sel ? S_S9_GNT : s9_hready ? S_S9_DATA : S_S9_CMD;
                          m2_s9_cmd_last = m2_s9_wt_sel ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m2_nxt_st[48:0] = S_S9_WAIT;
                  end
       endcase
  end
  S_S10_WAIT:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       case(1'b1)
         ~m2_s10_hld: begin
                          m2_nxt_st[48:0] = m2_s10_wt_sel ? S_S10_GNT : s10_hready ? S_S10_DATA : S_S10_CMD;
                          m2_s10_cmd_last = m2_s10_wt_sel ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m2_nxt_st[48:0] = S_S10_WAIT;
                  end
       endcase
  end
  S_S11_WAIT:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       case(1'b1)
         ~m2_s11_hld: begin
                          m2_nxt_st[48:0] = m2_s11_wt_sel ? S_S11_GNT : s11_hready ? S_S11_DATA : S_S11_CMD;
                          m2_s11_cmd_last = m2_s11_wt_sel ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m2_nxt_st[48:0] = S_S11_WAIT;
                  end
       endcase
  end
  S_S0_CMD: begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = s0_hready ? 1'b1 : 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       m2_nxt_st[48:0] = s0_hready  ? S_S0_DATA : S_S0_CMD;
  end
  S_S0_DATA:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b1;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       if(s0_hready)
         begin
           case(1'b1)
             m2_s0_sel: begin
                              m2_nxt_st[48:0] = S_S0_DATA;
                              m2_s0_cmd_cur = 1'b1;
                             end
             m2_s0_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S0_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s1_sel: begin
                              m2_nxt_st[48:0] = m2_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m2_latch_cmd = m2_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m2_s1_cmd_cur = m2_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m2_s1_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S1_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s2_sel: begin
                              m2_nxt_st[48:0] = m2_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m2_latch_cmd = m2_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m2_s2_cmd_cur = m2_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m2_s2_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S2_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s3_sel: begin
                              m2_nxt_st[48:0] = m2_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m2_latch_cmd = m2_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m2_s3_cmd_cur = m2_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m2_s3_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S3_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s4_sel: begin
                              m2_nxt_st[48:0] = m2_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m2_latch_cmd = m2_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m2_s4_cmd_cur = m2_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m2_s4_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S4_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s5_sel: begin
                              m2_nxt_st[48:0] = m2_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m2_latch_cmd = m2_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m2_s5_cmd_cur = m2_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m2_s5_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S5_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s6_sel: begin
                              m2_nxt_st[48:0] = m2_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m2_latch_cmd = m2_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m2_s6_cmd_cur = m2_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m2_s6_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S6_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s7_sel: begin
                              m2_nxt_st[48:0] = m2_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m2_latch_cmd = m2_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m2_s7_cmd_cur = m2_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m2_s7_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S7_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s8_sel: begin
                              m2_nxt_st[48:0] = m2_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m2_latch_cmd = m2_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m2_s8_cmd_cur = m2_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m2_s8_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S8_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s9_sel: begin
                              m2_nxt_st[48:0] = m2_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m2_latch_cmd = m2_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m2_s9_cmd_cur = m2_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m2_s9_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S9_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s10_sel: begin
                              m2_nxt_st[48:0] = m2_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m2_latch_cmd = m2_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m2_s10_cmd_cur = m2_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m2_s10_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S10_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s11_sel: begin
                              m2_nxt_st[48:0] = m2_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m2_latch_cmd = m2_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m2_s11_cmd_cur = m2_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m2_s11_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S11_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             default: begin
                             m2_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m2_nxt_st[48:0] = S_S0_DATA;
end
  S_S1_CMD: begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = s1_hready ? 1'b1 : 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       m2_nxt_st[48:0] = s1_hready  ? S_S1_DATA : S_S1_CMD;
  end
  S_S1_DATA:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b1;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       if(s1_hready)
         begin
           case(1'b1)
             m2_s0_sel: begin
                              m2_nxt_st[48:0] = m2_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m2_latch_cmd = m2_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m2_s0_cmd_cur = m2_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m2_s0_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S0_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s1_sel: begin
                              m2_nxt_st[48:0] = S_S1_DATA;
                              m2_s1_cmd_cur = 1'b1;
                             end
             m2_s1_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S1_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s2_sel: begin
                              m2_nxt_st[48:0] = m2_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m2_latch_cmd = m2_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m2_s2_cmd_cur = m2_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m2_s2_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S2_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s3_sel: begin
                              m2_nxt_st[48:0] = m2_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m2_latch_cmd = m2_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m2_s3_cmd_cur = m2_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m2_s3_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S3_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s4_sel: begin
                              m2_nxt_st[48:0] = m2_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m2_latch_cmd = m2_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m2_s4_cmd_cur = m2_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m2_s4_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S4_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s5_sel: begin
                              m2_nxt_st[48:0] = m2_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m2_latch_cmd = m2_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m2_s5_cmd_cur = m2_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m2_s5_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S5_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s6_sel: begin
                              m2_nxt_st[48:0] = m2_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m2_latch_cmd = m2_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m2_s6_cmd_cur = m2_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m2_s6_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S6_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s7_sel: begin
                              m2_nxt_st[48:0] = m2_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m2_latch_cmd = m2_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m2_s7_cmd_cur = m2_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m2_s7_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S7_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s8_sel: begin
                              m2_nxt_st[48:0] = m2_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m2_latch_cmd = m2_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m2_s8_cmd_cur = m2_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m2_s8_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S8_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s9_sel: begin
                              m2_nxt_st[48:0] = m2_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m2_latch_cmd = m2_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m2_s9_cmd_cur = m2_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m2_s9_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S9_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s10_sel: begin
                              m2_nxt_st[48:0] = m2_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m2_latch_cmd = m2_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m2_s10_cmd_cur = m2_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m2_s10_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S10_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s11_sel: begin
                              m2_nxt_st[48:0] = m2_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m2_latch_cmd = m2_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m2_s11_cmd_cur = m2_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m2_s11_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S11_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             default: begin
                             m2_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m2_nxt_st[48:0] = S_S1_DATA;
end
  S_S2_CMD: begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = s2_hready ? 1'b1 : 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       m2_nxt_st[48:0] = s2_hready  ? S_S2_DATA : S_S2_CMD;
  end
  S_S2_DATA:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b1;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       if(s2_hready)
         begin
           case(1'b1)
             m2_s0_sel: begin
                              m2_nxt_st[48:0] = m2_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m2_latch_cmd = m2_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m2_s0_cmd_cur = m2_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m2_s0_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S0_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s1_sel: begin
                              m2_nxt_st[48:0] = m2_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m2_latch_cmd = m2_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m2_s1_cmd_cur = m2_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m2_s1_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S1_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s2_sel: begin
                              m2_nxt_st[48:0] = S_S2_DATA;
                              m2_s2_cmd_cur = 1'b1;
                             end
             m2_s2_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S2_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s3_sel: begin
                              m2_nxt_st[48:0] = m2_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m2_latch_cmd = m2_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m2_s3_cmd_cur = m2_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m2_s3_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S3_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s4_sel: begin
                              m2_nxt_st[48:0] = m2_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m2_latch_cmd = m2_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m2_s4_cmd_cur = m2_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m2_s4_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S4_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s5_sel: begin
                              m2_nxt_st[48:0] = m2_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m2_latch_cmd = m2_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m2_s5_cmd_cur = m2_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m2_s5_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S5_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s6_sel: begin
                              m2_nxt_st[48:0] = m2_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m2_latch_cmd = m2_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m2_s6_cmd_cur = m2_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m2_s6_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S6_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s7_sel: begin
                              m2_nxt_st[48:0] = m2_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m2_latch_cmd = m2_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m2_s7_cmd_cur = m2_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m2_s7_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S7_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s8_sel: begin
                              m2_nxt_st[48:0] = m2_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m2_latch_cmd = m2_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m2_s8_cmd_cur = m2_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m2_s8_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S8_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s9_sel: begin
                              m2_nxt_st[48:0] = m2_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m2_latch_cmd = m2_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m2_s9_cmd_cur = m2_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m2_s9_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S9_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s10_sel: begin
                              m2_nxt_st[48:0] = m2_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m2_latch_cmd = m2_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m2_s10_cmd_cur = m2_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m2_s10_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S10_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s11_sel: begin
                              m2_nxt_st[48:0] = m2_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m2_latch_cmd = m2_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m2_s11_cmd_cur = m2_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m2_s11_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S11_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             default: begin
                             m2_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m2_nxt_st[48:0] = S_S2_DATA;
end
  S_S3_CMD: begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = s3_hready ? 1'b1 : 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       m2_nxt_st[48:0] = s3_hready  ? S_S3_DATA : S_S3_CMD;
  end
  S_S3_DATA:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b1;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       if(s3_hready)
         begin
           case(1'b1)
             m2_s0_sel: begin
                              m2_nxt_st[48:0] = m2_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m2_latch_cmd = m2_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m2_s0_cmd_cur = m2_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m2_s0_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S0_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s1_sel: begin
                              m2_nxt_st[48:0] = m2_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m2_latch_cmd = m2_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m2_s1_cmd_cur = m2_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m2_s1_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S1_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s2_sel: begin
                              m2_nxt_st[48:0] = m2_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m2_latch_cmd = m2_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m2_s2_cmd_cur = m2_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m2_s2_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S2_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s3_sel: begin
                              m2_nxt_st[48:0] = S_S3_DATA;
                              m2_s3_cmd_cur = 1'b1;
                             end
             m2_s3_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S3_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s4_sel: begin
                              m2_nxt_st[48:0] = m2_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m2_latch_cmd = m2_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m2_s4_cmd_cur = m2_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m2_s4_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S4_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s5_sel: begin
                              m2_nxt_st[48:0] = m2_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m2_latch_cmd = m2_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m2_s5_cmd_cur = m2_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m2_s5_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S5_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s6_sel: begin
                              m2_nxt_st[48:0] = m2_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m2_latch_cmd = m2_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m2_s6_cmd_cur = m2_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m2_s6_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S6_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s7_sel: begin
                              m2_nxt_st[48:0] = m2_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m2_latch_cmd = m2_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m2_s7_cmd_cur = m2_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m2_s7_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S7_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s8_sel: begin
                              m2_nxt_st[48:0] = m2_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m2_latch_cmd = m2_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m2_s8_cmd_cur = m2_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m2_s8_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S8_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s9_sel: begin
                              m2_nxt_st[48:0] = m2_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m2_latch_cmd = m2_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m2_s9_cmd_cur = m2_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m2_s9_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S9_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s10_sel: begin
                              m2_nxt_st[48:0] = m2_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m2_latch_cmd = m2_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m2_s10_cmd_cur = m2_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m2_s10_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S10_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s11_sel: begin
                              m2_nxt_st[48:0] = m2_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m2_latch_cmd = m2_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m2_s11_cmd_cur = m2_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m2_s11_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S11_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             default: begin
                             m2_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m2_nxt_st[48:0] = S_S3_DATA;
end
  S_S4_CMD: begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = s4_hready ? 1'b1 : 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       m2_nxt_st[48:0] = s4_hready  ? S_S4_DATA : S_S4_CMD;
  end
  S_S4_DATA:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b1;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       if(s4_hready)
         begin
           case(1'b1)
             m2_s0_sel: begin
                              m2_nxt_st[48:0] = m2_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m2_latch_cmd = m2_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m2_s0_cmd_cur = m2_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m2_s0_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S0_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s1_sel: begin
                              m2_nxt_st[48:0] = m2_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m2_latch_cmd = m2_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m2_s1_cmd_cur = m2_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m2_s1_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S1_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s2_sel: begin
                              m2_nxt_st[48:0] = m2_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m2_latch_cmd = m2_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m2_s2_cmd_cur = m2_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m2_s2_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S2_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s3_sel: begin
                              m2_nxt_st[48:0] = m2_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m2_latch_cmd = m2_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m2_s3_cmd_cur = m2_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m2_s3_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S3_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s4_sel: begin
                              m2_nxt_st[48:0] = S_S4_DATA;
                              m2_s4_cmd_cur = 1'b1;
                             end
             m2_s4_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S4_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s5_sel: begin
                              m2_nxt_st[48:0] = m2_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m2_latch_cmd = m2_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m2_s5_cmd_cur = m2_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m2_s5_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S5_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s6_sel: begin
                              m2_nxt_st[48:0] = m2_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m2_latch_cmd = m2_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m2_s6_cmd_cur = m2_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m2_s6_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S6_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s7_sel: begin
                              m2_nxt_st[48:0] = m2_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m2_latch_cmd = m2_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m2_s7_cmd_cur = m2_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m2_s7_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S7_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s8_sel: begin
                              m2_nxt_st[48:0] = m2_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m2_latch_cmd = m2_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m2_s8_cmd_cur = m2_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m2_s8_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S8_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s9_sel: begin
                              m2_nxt_st[48:0] = m2_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m2_latch_cmd = m2_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m2_s9_cmd_cur = m2_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m2_s9_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S9_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s10_sel: begin
                              m2_nxt_st[48:0] = m2_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m2_latch_cmd = m2_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m2_s10_cmd_cur = m2_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m2_s10_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S10_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s11_sel: begin
                              m2_nxt_st[48:0] = m2_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m2_latch_cmd = m2_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m2_s11_cmd_cur = m2_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m2_s11_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S11_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             default: begin
                             m2_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m2_nxt_st[48:0] = S_S4_DATA;
end
  S_S5_CMD: begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = s5_hready ? 1'b1 : 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       m2_nxt_st[48:0] = s5_hready  ? S_S5_DATA : S_S5_CMD;
  end
  S_S5_DATA:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b1;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       if(s5_hready)
         begin
           case(1'b1)
             m2_s0_sel: begin
                              m2_nxt_st[48:0] = m2_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m2_latch_cmd = m2_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m2_s0_cmd_cur = m2_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m2_s0_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S0_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s1_sel: begin
                              m2_nxt_st[48:0] = m2_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m2_latch_cmd = m2_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m2_s1_cmd_cur = m2_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m2_s1_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S1_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s2_sel: begin
                              m2_nxt_st[48:0] = m2_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m2_latch_cmd = m2_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m2_s2_cmd_cur = m2_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m2_s2_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S2_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s3_sel: begin
                              m2_nxt_st[48:0] = m2_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m2_latch_cmd = m2_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m2_s3_cmd_cur = m2_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m2_s3_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S3_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s4_sel: begin
                              m2_nxt_st[48:0] = m2_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m2_latch_cmd = m2_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m2_s4_cmd_cur = m2_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m2_s4_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S4_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s5_sel: begin
                              m2_nxt_st[48:0] = S_S5_DATA;
                              m2_s5_cmd_cur = 1'b1;
                             end
             m2_s5_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S5_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s6_sel: begin
                              m2_nxt_st[48:0] = m2_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m2_latch_cmd = m2_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m2_s6_cmd_cur = m2_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m2_s6_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S6_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s7_sel: begin
                              m2_nxt_st[48:0] = m2_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m2_latch_cmd = m2_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m2_s7_cmd_cur = m2_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m2_s7_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S7_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s8_sel: begin
                              m2_nxt_st[48:0] = m2_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m2_latch_cmd = m2_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m2_s8_cmd_cur = m2_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m2_s8_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S8_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s9_sel: begin
                              m2_nxt_st[48:0] = m2_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m2_latch_cmd = m2_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m2_s9_cmd_cur = m2_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m2_s9_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S9_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s10_sel: begin
                              m2_nxt_st[48:0] = m2_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m2_latch_cmd = m2_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m2_s10_cmd_cur = m2_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m2_s10_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S10_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s11_sel: begin
                              m2_nxt_st[48:0] = m2_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m2_latch_cmd = m2_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m2_s11_cmd_cur = m2_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m2_s11_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S11_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             default: begin
                             m2_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m2_nxt_st[48:0] = S_S5_DATA;
end
  S_S6_CMD: begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = s6_hready ? 1'b1 : 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       m2_nxt_st[48:0] = s6_hready  ? S_S6_DATA : S_S6_CMD;
  end
  S_S6_DATA:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b1;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       if(s6_hready)
         begin
           case(1'b1)
             m2_s0_sel: begin
                              m2_nxt_st[48:0] = m2_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m2_latch_cmd = m2_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m2_s0_cmd_cur = m2_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m2_s0_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S0_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s1_sel: begin
                              m2_nxt_st[48:0] = m2_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m2_latch_cmd = m2_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m2_s1_cmd_cur = m2_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m2_s1_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S1_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s2_sel: begin
                              m2_nxt_st[48:0] = m2_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m2_latch_cmd = m2_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m2_s2_cmd_cur = m2_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m2_s2_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S2_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s3_sel: begin
                              m2_nxt_st[48:0] = m2_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m2_latch_cmd = m2_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m2_s3_cmd_cur = m2_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m2_s3_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S3_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s4_sel: begin
                              m2_nxt_st[48:0] = m2_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m2_latch_cmd = m2_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m2_s4_cmd_cur = m2_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m2_s4_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S4_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s5_sel: begin
                              m2_nxt_st[48:0] = m2_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m2_latch_cmd = m2_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m2_s5_cmd_cur = m2_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m2_s5_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S5_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s6_sel: begin
                              m2_nxt_st[48:0] = S_S6_DATA;
                              m2_s6_cmd_cur = 1'b1;
                             end
             m2_s6_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S6_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s7_sel: begin
                              m2_nxt_st[48:0] = m2_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m2_latch_cmd = m2_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m2_s7_cmd_cur = m2_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m2_s7_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S7_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s8_sel: begin
                              m2_nxt_st[48:0] = m2_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m2_latch_cmd = m2_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m2_s8_cmd_cur = m2_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m2_s8_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S8_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s9_sel: begin
                              m2_nxt_st[48:0] = m2_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m2_latch_cmd = m2_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m2_s9_cmd_cur = m2_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m2_s9_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S9_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s10_sel: begin
                              m2_nxt_st[48:0] = m2_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m2_latch_cmd = m2_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m2_s10_cmd_cur = m2_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m2_s10_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S10_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s11_sel: begin
                              m2_nxt_st[48:0] = m2_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m2_latch_cmd = m2_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m2_s11_cmd_cur = m2_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m2_s11_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S11_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             default: begin
                             m2_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m2_nxt_st[48:0] = S_S6_DATA;
end
  S_S7_CMD: begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = s7_hready ? 1'b1 : 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       m2_nxt_st[48:0] = s7_hready  ? S_S7_DATA : S_S7_CMD;
  end
  S_S7_DATA:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b1;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       if(s7_hready)
         begin
           case(1'b1)
             m2_s0_sel: begin
                              m2_nxt_st[48:0] = m2_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m2_latch_cmd = m2_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m2_s0_cmd_cur = m2_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m2_s0_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S0_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s1_sel: begin
                              m2_nxt_st[48:0] = m2_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m2_latch_cmd = m2_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m2_s1_cmd_cur = m2_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m2_s1_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S1_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s2_sel: begin
                              m2_nxt_st[48:0] = m2_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m2_latch_cmd = m2_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m2_s2_cmd_cur = m2_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m2_s2_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S2_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s3_sel: begin
                              m2_nxt_st[48:0] = m2_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m2_latch_cmd = m2_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m2_s3_cmd_cur = m2_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m2_s3_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S3_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s4_sel: begin
                              m2_nxt_st[48:0] = m2_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m2_latch_cmd = m2_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m2_s4_cmd_cur = m2_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m2_s4_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S4_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s5_sel: begin
                              m2_nxt_st[48:0] = m2_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m2_latch_cmd = m2_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m2_s5_cmd_cur = m2_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m2_s5_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S5_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s6_sel: begin
                              m2_nxt_st[48:0] = m2_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m2_latch_cmd = m2_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m2_s6_cmd_cur = m2_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m2_s6_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S6_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s7_sel: begin
                              m2_nxt_st[48:0] = S_S7_DATA;
                              m2_s7_cmd_cur = 1'b1;
                             end
             m2_s7_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S7_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s8_sel: begin
                              m2_nxt_st[48:0] = m2_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m2_latch_cmd = m2_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m2_s8_cmd_cur = m2_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m2_s8_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S8_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s9_sel: begin
                              m2_nxt_st[48:0] = m2_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m2_latch_cmd = m2_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m2_s9_cmd_cur = m2_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m2_s9_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S9_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s10_sel: begin
                              m2_nxt_st[48:0] = m2_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m2_latch_cmd = m2_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m2_s10_cmd_cur = m2_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m2_s10_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S10_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s11_sel: begin
                              m2_nxt_st[48:0] = m2_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m2_latch_cmd = m2_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m2_s11_cmd_cur = m2_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m2_s11_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S11_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             default: begin
                             m2_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m2_nxt_st[48:0] = S_S7_DATA;
end
  S_S8_CMD: begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = s8_hready ? 1'b1 : 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       m2_nxt_st[48:0] = s8_hready  ? S_S8_DATA : S_S8_CMD;
  end
  S_S8_DATA:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b1;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       if(s8_hready)
         begin
           case(1'b1)
             m2_s0_sel: begin
                              m2_nxt_st[48:0] = m2_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m2_latch_cmd = m2_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m2_s0_cmd_cur = m2_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m2_s0_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S0_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s1_sel: begin
                              m2_nxt_st[48:0] = m2_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m2_latch_cmd = m2_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m2_s1_cmd_cur = m2_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m2_s1_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S1_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s2_sel: begin
                              m2_nxt_st[48:0] = m2_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m2_latch_cmd = m2_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m2_s2_cmd_cur = m2_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m2_s2_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S2_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s3_sel: begin
                              m2_nxt_st[48:0] = m2_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m2_latch_cmd = m2_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m2_s3_cmd_cur = m2_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m2_s3_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S3_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s4_sel: begin
                              m2_nxt_st[48:0] = m2_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m2_latch_cmd = m2_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m2_s4_cmd_cur = m2_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m2_s4_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S4_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s5_sel: begin
                              m2_nxt_st[48:0] = m2_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m2_latch_cmd = m2_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m2_s5_cmd_cur = m2_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m2_s5_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S5_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s6_sel: begin
                              m2_nxt_st[48:0] = m2_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m2_latch_cmd = m2_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m2_s6_cmd_cur = m2_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m2_s6_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S6_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s7_sel: begin
                              m2_nxt_st[48:0] = m2_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m2_latch_cmd = m2_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m2_s7_cmd_cur = m2_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m2_s7_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S7_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s8_sel: begin
                              m2_nxt_st[48:0] = S_S8_DATA;
                              m2_s8_cmd_cur = 1'b1;
                             end
             m2_s8_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S8_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s9_sel: begin
                              m2_nxt_st[48:0] = m2_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m2_latch_cmd = m2_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m2_s9_cmd_cur = m2_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m2_s9_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S9_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s10_sel: begin
                              m2_nxt_st[48:0] = m2_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m2_latch_cmd = m2_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m2_s10_cmd_cur = m2_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m2_s10_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S10_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s11_sel: begin
                              m2_nxt_st[48:0] = m2_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m2_latch_cmd = m2_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m2_s11_cmd_cur = m2_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m2_s11_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S11_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             default: begin
                             m2_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m2_nxt_st[48:0] = S_S8_DATA;
end
  S_S9_CMD: begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = s9_hready ? 1'b1 : 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       m2_nxt_st[48:0] = s9_hready  ? S_S9_DATA : S_S9_CMD;
  end
  S_S9_DATA:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b1;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       if(s9_hready)
         begin
           case(1'b1)
             m2_s0_sel: begin
                              m2_nxt_st[48:0] = m2_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m2_latch_cmd = m2_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m2_s0_cmd_cur = m2_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m2_s0_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S0_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s1_sel: begin
                              m2_nxt_st[48:0] = m2_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m2_latch_cmd = m2_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m2_s1_cmd_cur = m2_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m2_s1_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S1_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s2_sel: begin
                              m2_nxt_st[48:0] = m2_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m2_latch_cmd = m2_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m2_s2_cmd_cur = m2_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m2_s2_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S2_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s3_sel: begin
                              m2_nxt_st[48:0] = m2_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m2_latch_cmd = m2_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m2_s3_cmd_cur = m2_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m2_s3_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S3_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s4_sel: begin
                              m2_nxt_st[48:0] = m2_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m2_latch_cmd = m2_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m2_s4_cmd_cur = m2_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m2_s4_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S4_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s5_sel: begin
                              m2_nxt_st[48:0] = m2_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m2_latch_cmd = m2_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m2_s5_cmd_cur = m2_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m2_s5_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S5_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s6_sel: begin
                              m2_nxt_st[48:0] = m2_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m2_latch_cmd = m2_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m2_s6_cmd_cur = m2_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m2_s6_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S6_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s7_sel: begin
                              m2_nxt_st[48:0] = m2_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m2_latch_cmd = m2_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m2_s7_cmd_cur = m2_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m2_s7_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S7_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s8_sel: begin
                              m2_nxt_st[48:0] = m2_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m2_latch_cmd = m2_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m2_s8_cmd_cur = m2_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m2_s8_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S8_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s9_sel: begin
                              m2_nxt_st[48:0] = S_S9_DATA;
                              m2_s9_cmd_cur = 1'b1;
                             end
             m2_s9_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S9_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s10_sel: begin
                              m2_nxt_st[48:0] = m2_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m2_latch_cmd = m2_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m2_s10_cmd_cur = m2_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m2_s10_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S10_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s11_sel: begin
                              m2_nxt_st[48:0] = m2_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m2_latch_cmd = m2_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m2_s11_cmd_cur = m2_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m2_s11_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S11_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             default: begin
                             m2_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m2_nxt_st[48:0] = S_S9_DATA;
end
  S_S10_CMD: begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = s10_hready ? 1'b1 : 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       m2_nxt_st[48:0] = s10_hready  ? S_S10_DATA : S_S10_CMD;
  end
  S_S10_DATA:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b1;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       if(s10_hready)
         begin
           case(1'b1)
             m2_s0_sel: begin
                              m2_nxt_st[48:0] = m2_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m2_latch_cmd = m2_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m2_s0_cmd_cur = m2_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m2_s0_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S0_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s1_sel: begin
                              m2_nxt_st[48:0] = m2_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m2_latch_cmd = m2_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m2_s1_cmd_cur = m2_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m2_s1_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S1_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s2_sel: begin
                              m2_nxt_st[48:0] = m2_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m2_latch_cmd = m2_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m2_s2_cmd_cur = m2_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m2_s2_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S2_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s3_sel: begin
                              m2_nxt_st[48:0] = m2_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m2_latch_cmd = m2_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m2_s3_cmd_cur = m2_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m2_s3_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S3_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s4_sel: begin
                              m2_nxt_st[48:0] = m2_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m2_latch_cmd = m2_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m2_s4_cmd_cur = m2_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m2_s4_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S4_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s5_sel: begin
                              m2_nxt_st[48:0] = m2_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m2_latch_cmd = m2_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m2_s5_cmd_cur = m2_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m2_s5_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S5_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s6_sel: begin
                              m2_nxt_st[48:0] = m2_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m2_latch_cmd = m2_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m2_s6_cmd_cur = m2_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m2_s6_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S6_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s7_sel: begin
                              m2_nxt_st[48:0] = m2_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m2_latch_cmd = m2_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m2_s7_cmd_cur = m2_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m2_s7_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S7_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s8_sel: begin
                              m2_nxt_st[48:0] = m2_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m2_latch_cmd = m2_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m2_s8_cmd_cur = m2_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m2_s8_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S8_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s9_sel: begin
                              m2_nxt_st[48:0] = m2_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m2_latch_cmd = m2_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m2_s9_cmd_cur = m2_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m2_s9_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S9_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s10_sel: begin
                              m2_nxt_st[48:0] = S_S10_DATA;
                              m2_s10_cmd_cur = 1'b1;
                             end
             m2_s10_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S10_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s11_sel: begin
                              m2_nxt_st[48:0] = m2_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m2_latch_cmd = m2_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m2_s11_cmd_cur = m2_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m2_s11_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S11_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             default: begin
                             m2_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m2_nxt_st[48:0] = S_S10_DATA;
end
  S_S11_CMD: begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = s11_hready ? 1'b1 : 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b0;
       m2_nxt_st[48:0] = s11_hready  ? S_S11_DATA : S_S11_CMD;
  end
  S_S11_DATA:begin
       m2_latch_cmd = 1'b0;
       m2_s0_cmd_last = 1'b0;
       m2_s0_cmd_cur = 1'b0;
       m2_s0_data = 1'b0;
       m2_s1_cmd_last = 1'b0;
       m2_s1_cmd_cur = 1'b0;
       m2_s1_data = 1'b0;
       m2_s2_cmd_last = 1'b0;
       m2_s2_cmd_cur = 1'b0;
       m2_s2_data = 1'b0;
       m2_s3_cmd_last = 1'b0;
       m2_s3_cmd_cur = 1'b0;
       m2_s3_data = 1'b0;
       m2_s4_cmd_last = 1'b0;
       m2_s4_cmd_cur = 1'b0;
       m2_s4_data = 1'b0;
       m2_s5_cmd_last = 1'b0;
       m2_s5_cmd_cur = 1'b0;
       m2_s5_data = 1'b0;
       m2_s6_cmd_last = 1'b0;
       m2_s6_cmd_cur = 1'b0;
       m2_s6_data = 1'b0;
       m2_s7_cmd_last = 1'b0;
       m2_s7_cmd_cur = 1'b0;
       m2_s7_data = 1'b0;
       m2_s8_cmd_last = 1'b0;
       m2_s8_cmd_cur = 1'b0;
       m2_s8_data = 1'b0;
       m2_s9_cmd_last = 1'b0;
       m2_s9_cmd_cur = 1'b0;
       m2_s9_data = 1'b0;
       m2_s10_cmd_last = 1'b0;
       m2_s10_cmd_cur = 1'b0;
       m2_s10_data = 1'b0;
       m2_s11_cmd_last = 1'b0;
       m2_s11_cmd_cur = 1'b0;
       m2_s11_data = 1'b1;
       if(s11_hready)
         begin
           case(1'b1)
             m2_s0_sel: begin
                              m2_nxt_st[48:0] = m2_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m2_latch_cmd = m2_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m2_s0_cmd_cur = m2_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m2_s0_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S0_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s1_sel: begin
                              m2_nxt_st[48:0] = m2_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m2_latch_cmd = m2_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m2_s1_cmd_cur = m2_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m2_s1_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S1_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s2_sel: begin
                              m2_nxt_st[48:0] = m2_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m2_latch_cmd = m2_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m2_s2_cmd_cur = m2_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m2_s2_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S2_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s3_sel: begin
                              m2_nxt_st[48:0] = m2_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m2_latch_cmd = m2_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m2_s3_cmd_cur = m2_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m2_s3_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S3_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s4_sel: begin
                              m2_nxt_st[48:0] = m2_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m2_latch_cmd = m2_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m2_s4_cmd_cur = m2_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m2_s4_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S4_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s5_sel: begin
                              m2_nxt_st[48:0] = m2_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m2_latch_cmd = m2_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m2_s5_cmd_cur = m2_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m2_s5_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S5_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s6_sel: begin
                              m2_nxt_st[48:0] = m2_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m2_latch_cmd = m2_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m2_s6_cmd_cur = m2_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m2_s6_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S6_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s7_sel: begin
                              m2_nxt_st[48:0] = m2_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m2_latch_cmd = m2_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m2_s7_cmd_cur = m2_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m2_s7_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S7_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s8_sel: begin
                              m2_nxt_st[48:0] = m2_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m2_latch_cmd = m2_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m2_s8_cmd_cur = m2_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m2_s8_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S8_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s9_sel: begin
                              m2_nxt_st[48:0] = m2_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m2_latch_cmd = m2_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m2_s9_cmd_cur = m2_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m2_s9_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S9_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s10_sel: begin
                              m2_nxt_st[48:0] = m2_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m2_latch_cmd = m2_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m2_s10_cmd_cur = m2_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m2_s10_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S10_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             m2_s11_sel: begin
                              m2_nxt_st[48:0] = S_S11_DATA;
                              m2_s11_cmd_cur = 1'b1;
                             end
             m2_s11_wt_sel: begin
                                 m2_nxt_st[48:0] = S_S11_GNT;
                                 m2_latch_cmd = 1'b1;
                               end
             default: begin
                             m2_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m2_nxt_st[48:0] = S_S11_DATA;
end
  default: begin
             m2_latch_cmd = 1'b0;
             m2_s0_cmd_last = 1'b0;
             m2_s0_cmd_cur = 1'b0;
             m2_s0_data = 1'b0;
             m2_s1_cmd_last = 1'b0;
             m2_s1_cmd_cur = 1'b0;
             m2_s1_data = 1'b0;
             m2_s2_cmd_last = 1'b0;
             m2_s2_cmd_cur = 1'b0;
             m2_s2_data = 1'b0;
             m2_s3_cmd_last = 1'b0;
             m2_s3_cmd_cur = 1'b0;
             m2_s3_data = 1'b0;
             m2_s4_cmd_last = 1'b0;
             m2_s4_cmd_cur = 1'b0;
             m2_s4_data = 1'b0;
             m2_s5_cmd_last = 1'b0;
             m2_s5_cmd_cur = 1'b0;
             m2_s5_data = 1'b0;
             m2_s6_cmd_last = 1'b0;
             m2_s6_cmd_cur = 1'b0;
             m2_s6_data = 1'b0;
             m2_s7_cmd_last = 1'b0;
             m2_s7_cmd_cur = 1'b0;
             m2_s7_data = 1'b0;
             m2_s8_cmd_last = 1'b0;
             m2_s8_cmd_cur = 1'b0;
             m2_s8_data = 1'b0;
             m2_s9_cmd_last = 1'b0;
             m2_s9_cmd_cur = 1'b0;
             m2_s9_data = 1'b0;
             m2_s10_cmd_last = 1'b0;
             m2_s10_cmd_cur = 1'b0;
             m2_s10_data = 1'b0;
             m2_s11_cmd_last = 1'b0;
             m2_s11_cmd_cur = 1'b0;
             m2_s11_data = 1'b0;
             m2_nxt_st[48:0] = S_IDLE;
  end
endcase
end
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
       m3_cur_st[48:0] <= S_IDLE;
    else
       m3_cur_st[48:0] <= m3_nxt_st[48:0];
  end
always @ (*)
begin
case(m3_cur_st[48:0])
  S_IDLE:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       case(1'b1)
         m3_s0_sel: begin
                          m3_nxt_st[48:0] = m3_s0_hld ? S_S0_WAIT : (s0_hready ? S_S0_DATA : S_S0_CMD);
                          m3_latch_cmd = m3_s0_hld ? 1'b1 : (s0_hready ? 1'b0 : 1'b1);
                          m3_s0_cmd_cur = m3_s0_hld ? 1'b0 : (s0_hready ? 1'b1 : 1'b0);
                        end
         m3_s0_wt_sel: begin
                             m3_nxt_st[48:0] = S_S0_GNT;
                             m3_latch_cmd = 1'b1;
                           end
         m3_s1_sel: begin
                          m3_nxt_st[48:0] = m3_s1_hld ? S_S1_WAIT : (s1_hready ? S_S1_DATA : S_S1_CMD);
                          m3_latch_cmd = m3_s1_hld ? 1'b1 : (s1_hready ? 1'b0 : 1'b1);
                          m3_s1_cmd_cur = m3_s1_hld ? 1'b0 : (s1_hready ? 1'b1 : 1'b0);
                        end
         m3_s1_wt_sel: begin
                             m3_nxt_st[48:0] = S_S1_GNT;
                             m3_latch_cmd = 1'b1;
                           end
         m3_s2_sel: begin
                          m3_nxt_st[48:0] = m3_s2_hld ? S_S2_WAIT : (s2_hready ? S_S2_DATA : S_S2_CMD);
                          m3_latch_cmd = m3_s2_hld ? 1'b1 : (s2_hready ? 1'b0 : 1'b1);
                          m3_s2_cmd_cur = m3_s2_hld ? 1'b0 : (s2_hready ? 1'b1 : 1'b0);
                        end
         m3_s2_wt_sel: begin
                             m3_nxt_st[48:0] = S_S2_GNT;
                             m3_latch_cmd = 1'b1;
                           end
         m3_s3_sel: begin
                          m3_nxt_st[48:0] = m3_s3_hld ? S_S3_WAIT : (s3_hready ? S_S3_DATA : S_S3_CMD);
                          m3_latch_cmd = m3_s3_hld ? 1'b1 : (s3_hready ? 1'b0 : 1'b1);
                          m3_s3_cmd_cur = m3_s3_hld ? 1'b0 : (s3_hready ? 1'b1 : 1'b0);
                        end
         m3_s3_wt_sel: begin
                             m3_nxt_st[48:0] = S_S3_GNT;
                             m3_latch_cmd = 1'b1;
                           end
         m3_s4_sel: begin
                          m3_nxt_st[48:0] = m3_s4_hld ? S_S4_WAIT : (s4_hready ? S_S4_DATA : S_S4_CMD);
                          m3_latch_cmd = m3_s4_hld ? 1'b1 : (s4_hready ? 1'b0 : 1'b1);
                          m3_s4_cmd_cur = m3_s4_hld ? 1'b0 : (s4_hready ? 1'b1 : 1'b0);
                        end
         m3_s4_wt_sel: begin
                             m3_nxt_st[48:0] = S_S4_GNT;
                             m3_latch_cmd = 1'b1;
                           end
         m3_s5_sel: begin
                          m3_nxt_st[48:0] = m3_s5_hld ? S_S5_WAIT : (s5_hready ? S_S5_DATA : S_S5_CMD);
                          m3_latch_cmd = m3_s5_hld ? 1'b1 : (s5_hready ? 1'b0 : 1'b1);
                          m3_s5_cmd_cur = m3_s5_hld ? 1'b0 : (s5_hready ? 1'b1 : 1'b0);
                        end
         m3_s5_wt_sel: begin
                             m3_nxt_st[48:0] = S_S5_GNT;
                             m3_latch_cmd = 1'b1;
                           end
         m3_s6_sel: begin
                          m3_nxt_st[48:0] = m3_s6_hld ? S_S6_WAIT : (s6_hready ? S_S6_DATA : S_S6_CMD);
                          m3_latch_cmd = m3_s6_hld ? 1'b1 : (s6_hready ? 1'b0 : 1'b1);
                          m3_s6_cmd_cur = m3_s6_hld ? 1'b0 : (s6_hready ? 1'b1 : 1'b0);
                        end
         m3_s6_wt_sel: begin
                             m3_nxt_st[48:0] = S_S6_GNT;
                             m3_latch_cmd = 1'b1;
                           end
         m3_s7_sel: begin
                          m3_nxt_st[48:0] = m3_s7_hld ? S_S7_WAIT : (s7_hready ? S_S7_DATA : S_S7_CMD);
                          m3_latch_cmd = m3_s7_hld ? 1'b1 : (s7_hready ? 1'b0 : 1'b1);
                          m3_s7_cmd_cur = m3_s7_hld ? 1'b0 : (s7_hready ? 1'b1 : 1'b0);
                        end
         m3_s7_wt_sel: begin
                             m3_nxt_st[48:0] = S_S7_GNT;
                             m3_latch_cmd = 1'b1;
                           end
         m3_s8_sel: begin
                          m3_nxt_st[48:0] = m3_s8_hld ? S_S8_WAIT : (s8_hready ? S_S8_DATA : S_S8_CMD);
                          m3_latch_cmd = m3_s8_hld ? 1'b1 : (s8_hready ? 1'b0 : 1'b1);
                          m3_s8_cmd_cur = m3_s8_hld ? 1'b0 : (s8_hready ? 1'b1 : 1'b0);
                        end
         m3_s8_wt_sel: begin
                             m3_nxt_st[48:0] = S_S8_GNT;
                             m3_latch_cmd = 1'b1;
                           end
         m3_s9_sel: begin
                          m3_nxt_st[48:0] = m3_s9_hld ? S_S9_WAIT : (s9_hready ? S_S9_DATA : S_S9_CMD);
                          m3_latch_cmd = m3_s9_hld ? 1'b1 : (s9_hready ? 1'b0 : 1'b1);
                          m3_s9_cmd_cur = m3_s9_hld ? 1'b0 : (s9_hready ? 1'b1 : 1'b0);
                        end
         m3_s9_wt_sel: begin
                             m3_nxt_st[48:0] = S_S9_GNT;
                             m3_latch_cmd = 1'b1;
                           end
         m3_s10_sel: begin
                          m3_nxt_st[48:0] = m3_s10_hld ? S_S10_WAIT : (s10_hready ? S_S10_DATA : S_S10_CMD);
                          m3_latch_cmd = m3_s10_hld ? 1'b1 : (s10_hready ? 1'b0 : 1'b1);
                          m3_s10_cmd_cur = m3_s10_hld ? 1'b0 : (s10_hready ? 1'b1 : 1'b0);
                        end
         m3_s10_wt_sel: begin
                             m3_nxt_st[48:0] = S_S10_GNT;
                             m3_latch_cmd = 1'b1;
                           end
         m3_s11_sel: begin
                          m3_nxt_st[48:0] = m3_s11_hld ? S_S11_WAIT : (s11_hready ? S_S11_DATA : S_S11_CMD);
                          m3_latch_cmd = m3_s11_hld ? 1'b1 : (s11_hready ? 1'b0 : 1'b1);
                          m3_s11_cmd_cur = m3_s11_hld ? 1'b0 : (s11_hready ? 1'b1 : 1'b0);
                        end
         m3_s11_wt_sel: begin
                             m3_nxt_st[48:0] = S_S11_GNT;
                             m3_latch_cmd = 1'b1;
                           end
         default: begin
                          m3_nxt_st[48:0] = S_IDLE;
                  end
       endcase
  end
  S_S0_GNT:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       case(1'b1)
         m3_s0_sel: begin
                          m3_nxt_st[48:0] = m3_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                          m3_s0_cmd_last = m3_s0_hld ? 1'b0 : (s0_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m3_nxt_st[48:0] = S_S0_GNT;
                  end
       endcase
  end
  S_S1_GNT:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       case(1'b1)
         m3_s1_sel: begin
                          m3_nxt_st[48:0] = m3_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                          m3_s1_cmd_last = m3_s1_hld ? 1'b0 : (s1_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m3_nxt_st[48:0] = S_S1_GNT;
                  end
       endcase
  end
  S_S2_GNT:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       case(1'b1)
         m3_s2_sel: begin
                          m3_nxt_st[48:0] = m3_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                          m3_s2_cmd_last = m3_s2_hld ? 1'b0 : (s2_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m3_nxt_st[48:0] = S_S2_GNT;
                  end
       endcase
  end
  S_S3_GNT:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       case(1'b1)
         m3_s3_sel: begin
                          m3_nxt_st[48:0] = m3_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                          m3_s3_cmd_last = m3_s3_hld ? 1'b0 : (s3_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m3_nxt_st[48:0] = S_S3_GNT;
                  end
       endcase
  end
  S_S4_GNT:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       case(1'b1)
         m3_s4_sel: begin
                          m3_nxt_st[48:0] = m3_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                          m3_s4_cmd_last = m3_s4_hld ? 1'b0 : (s4_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m3_nxt_st[48:0] = S_S4_GNT;
                  end
       endcase
  end
  S_S5_GNT:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       case(1'b1)
         m3_s5_sel: begin
                          m3_nxt_st[48:0] = m3_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                          m3_s5_cmd_last = m3_s5_hld ? 1'b0 : (s5_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m3_nxt_st[48:0] = S_S5_GNT;
                  end
       endcase
  end
  S_S6_GNT:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       case(1'b1)
         m3_s6_sel: begin
                          m3_nxt_st[48:0] = m3_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                          m3_s6_cmd_last = m3_s6_hld ? 1'b0 : (s6_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m3_nxt_st[48:0] = S_S6_GNT;
                  end
       endcase
  end
  S_S7_GNT:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       case(1'b1)
         m3_s7_sel: begin
                          m3_nxt_st[48:0] = m3_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                          m3_s7_cmd_last = m3_s7_hld ? 1'b0 : (s7_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m3_nxt_st[48:0] = S_S7_GNT;
                  end
       endcase
  end
  S_S8_GNT:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       case(1'b1)
         m3_s8_sel: begin
                          m3_nxt_st[48:0] = m3_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                          m3_s8_cmd_last = m3_s8_hld ? 1'b0 : (s8_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m3_nxt_st[48:0] = S_S8_GNT;
                  end
       endcase
  end
  S_S9_GNT:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       case(1'b1)
         m3_s9_sel: begin
                          m3_nxt_st[48:0] = m3_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                          m3_s9_cmd_last = m3_s9_hld ? 1'b0 : (s9_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m3_nxt_st[48:0] = S_S9_GNT;
                  end
       endcase
  end
  S_S10_GNT:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       case(1'b1)
         m3_s10_sel: begin
                          m3_nxt_st[48:0] = m3_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                          m3_s10_cmd_last = m3_s10_hld ? 1'b0 : (s10_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m3_nxt_st[48:0] = S_S10_GNT;
                  end
       endcase
  end
  S_S11_GNT:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       case(1'b1)
         m3_s11_sel: begin
                          m3_nxt_st[48:0] = m3_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                          m3_s11_cmd_last = m3_s11_hld ? 1'b0 : (s11_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m3_nxt_st[48:0] = S_S11_GNT;
                  end
       endcase
  end
  S_S0_WAIT:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       case(1'b1)
         ~m3_s0_hld: begin
                          m3_nxt_st[48:0] = m3_s0_wt_sel ? S_S0_GNT : s0_hready ? S_S0_DATA : S_S0_CMD;
                          m3_s0_cmd_last = m3_s0_wt_sel ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m3_nxt_st[48:0] = S_S0_WAIT;
                  end
       endcase
  end
  S_S1_WAIT:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       case(1'b1)
         ~m3_s1_hld: begin
                          m3_nxt_st[48:0] = m3_s1_wt_sel ? S_S1_GNT : s1_hready ? S_S1_DATA : S_S1_CMD;
                          m3_s1_cmd_last = m3_s1_wt_sel ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m3_nxt_st[48:0] = S_S1_WAIT;
                  end
       endcase
  end
  S_S2_WAIT:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       case(1'b1)
         ~m3_s2_hld: begin
                          m3_nxt_st[48:0] = m3_s2_wt_sel ? S_S2_GNT : s2_hready ? S_S2_DATA : S_S2_CMD;
                          m3_s2_cmd_last = m3_s2_wt_sel ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m3_nxt_st[48:0] = S_S2_WAIT;
                  end
       endcase
  end
  S_S3_WAIT:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       case(1'b1)
         ~m3_s3_hld: begin
                          m3_nxt_st[48:0] = m3_s3_wt_sel ? S_S3_GNT : s3_hready ? S_S3_DATA : S_S3_CMD;
                          m3_s3_cmd_last = m3_s3_wt_sel ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m3_nxt_st[48:0] = S_S3_WAIT;
                  end
       endcase
  end
  S_S4_WAIT:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       case(1'b1)
         ~m3_s4_hld: begin
                          m3_nxt_st[48:0] = m3_s4_wt_sel ? S_S4_GNT : s4_hready ? S_S4_DATA : S_S4_CMD;
                          m3_s4_cmd_last = m3_s4_wt_sel ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m3_nxt_st[48:0] = S_S4_WAIT;
                  end
       endcase
  end
  S_S5_WAIT:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       case(1'b1)
         ~m3_s5_hld: begin
                          m3_nxt_st[48:0] = m3_s5_wt_sel ? S_S5_GNT : s5_hready ? S_S5_DATA : S_S5_CMD;
                          m3_s5_cmd_last = m3_s5_wt_sel ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m3_nxt_st[48:0] = S_S5_WAIT;
                  end
       endcase
  end
  S_S6_WAIT:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       case(1'b1)
         ~m3_s6_hld: begin
                          m3_nxt_st[48:0] = m3_s6_wt_sel ? S_S6_GNT : s6_hready ? S_S6_DATA : S_S6_CMD;
                          m3_s6_cmd_last = m3_s6_wt_sel ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m3_nxt_st[48:0] = S_S6_WAIT;
                  end
       endcase
  end
  S_S7_WAIT:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       case(1'b1)
         ~m3_s7_hld: begin
                          m3_nxt_st[48:0] = m3_s7_wt_sel ? S_S7_GNT : s7_hready ? S_S7_DATA : S_S7_CMD;
                          m3_s7_cmd_last = m3_s7_wt_sel ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m3_nxt_st[48:0] = S_S7_WAIT;
                  end
       endcase
  end
  S_S8_WAIT:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       case(1'b1)
         ~m3_s8_hld: begin
                          m3_nxt_st[48:0] = m3_s8_wt_sel ? S_S8_GNT : s8_hready ? S_S8_DATA : S_S8_CMD;
                          m3_s8_cmd_last = m3_s8_wt_sel ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m3_nxt_st[48:0] = S_S8_WAIT;
                  end
       endcase
  end
  S_S9_WAIT:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       case(1'b1)
         ~m3_s9_hld: begin
                          m3_nxt_st[48:0] = m3_s9_wt_sel ? S_S9_GNT : s9_hready ? S_S9_DATA : S_S9_CMD;
                          m3_s9_cmd_last = m3_s9_wt_sel ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m3_nxt_st[48:0] = S_S9_WAIT;
                  end
       endcase
  end
  S_S10_WAIT:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       case(1'b1)
         ~m3_s10_hld: begin
                          m3_nxt_st[48:0] = m3_s10_wt_sel ? S_S10_GNT : s10_hready ? S_S10_DATA : S_S10_CMD;
                          m3_s10_cmd_last = m3_s10_wt_sel ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m3_nxt_st[48:0] = S_S10_WAIT;
                  end
       endcase
  end
  S_S11_WAIT:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       case(1'b1)
         ~m3_s11_hld: begin
                          m3_nxt_st[48:0] = m3_s11_wt_sel ? S_S11_GNT : s11_hready ? S_S11_DATA : S_S11_CMD;
                          m3_s11_cmd_last = m3_s11_wt_sel ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m3_nxt_st[48:0] = S_S11_WAIT;
                  end
       endcase
  end
  S_S0_CMD: begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = s0_hready ? 1'b1 : 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       m3_nxt_st[48:0] = s0_hready  ? S_S0_DATA : S_S0_CMD;
  end
  S_S0_DATA:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b1;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       if(s0_hready)
         begin
           case(1'b1)
             m3_s0_sel: begin
                              m3_nxt_st[48:0] = S_S0_DATA;
                              m3_s0_cmd_cur = 1'b1;
                             end
             m3_s0_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S0_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s1_sel: begin
                              m3_nxt_st[48:0] = m3_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m3_latch_cmd = m3_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m3_s1_cmd_cur = m3_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m3_s1_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S1_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s2_sel: begin
                              m3_nxt_st[48:0] = m3_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m3_latch_cmd = m3_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m3_s2_cmd_cur = m3_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m3_s2_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S2_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s3_sel: begin
                              m3_nxt_st[48:0] = m3_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m3_latch_cmd = m3_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m3_s3_cmd_cur = m3_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m3_s3_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S3_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s4_sel: begin
                              m3_nxt_st[48:0] = m3_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m3_latch_cmd = m3_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m3_s4_cmd_cur = m3_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m3_s4_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S4_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s5_sel: begin
                              m3_nxt_st[48:0] = m3_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m3_latch_cmd = m3_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m3_s5_cmd_cur = m3_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m3_s5_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S5_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s6_sel: begin
                              m3_nxt_st[48:0] = m3_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m3_latch_cmd = m3_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m3_s6_cmd_cur = m3_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m3_s6_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S6_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s7_sel: begin
                              m3_nxt_st[48:0] = m3_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m3_latch_cmd = m3_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m3_s7_cmd_cur = m3_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m3_s7_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S7_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s8_sel: begin
                              m3_nxt_st[48:0] = m3_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m3_latch_cmd = m3_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m3_s8_cmd_cur = m3_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m3_s8_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S8_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s9_sel: begin
                              m3_nxt_st[48:0] = m3_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m3_latch_cmd = m3_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m3_s9_cmd_cur = m3_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m3_s9_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S9_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s10_sel: begin
                              m3_nxt_st[48:0] = m3_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m3_latch_cmd = m3_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m3_s10_cmd_cur = m3_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m3_s10_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S10_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s11_sel: begin
                              m3_nxt_st[48:0] = m3_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m3_latch_cmd = m3_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m3_s11_cmd_cur = m3_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m3_s11_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S11_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             default: begin
                             m3_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m3_nxt_st[48:0] = S_S0_DATA;
end
  S_S1_CMD: begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = s1_hready ? 1'b1 : 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       m3_nxt_st[48:0] = s1_hready  ? S_S1_DATA : S_S1_CMD;
  end
  S_S1_DATA:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b1;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       if(s1_hready)
         begin
           case(1'b1)
             m3_s0_sel: begin
                              m3_nxt_st[48:0] = m3_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m3_latch_cmd = m3_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m3_s0_cmd_cur = m3_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m3_s0_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S0_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s1_sel: begin
                              m3_nxt_st[48:0] = S_S1_DATA;
                              m3_s1_cmd_cur = 1'b1;
                             end
             m3_s1_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S1_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s2_sel: begin
                              m3_nxt_st[48:0] = m3_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m3_latch_cmd = m3_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m3_s2_cmd_cur = m3_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m3_s2_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S2_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s3_sel: begin
                              m3_nxt_st[48:0] = m3_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m3_latch_cmd = m3_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m3_s3_cmd_cur = m3_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m3_s3_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S3_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s4_sel: begin
                              m3_nxt_st[48:0] = m3_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m3_latch_cmd = m3_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m3_s4_cmd_cur = m3_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m3_s4_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S4_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s5_sel: begin
                              m3_nxt_st[48:0] = m3_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m3_latch_cmd = m3_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m3_s5_cmd_cur = m3_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m3_s5_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S5_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s6_sel: begin
                              m3_nxt_st[48:0] = m3_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m3_latch_cmd = m3_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m3_s6_cmd_cur = m3_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m3_s6_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S6_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s7_sel: begin
                              m3_nxt_st[48:0] = m3_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m3_latch_cmd = m3_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m3_s7_cmd_cur = m3_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m3_s7_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S7_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s8_sel: begin
                              m3_nxt_st[48:0] = m3_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m3_latch_cmd = m3_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m3_s8_cmd_cur = m3_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m3_s8_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S8_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s9_sel: begin
                              m3_nxt_st[48:0] = m3_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m3_latch_cmd = m3_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m3_s9_cmd_cur = m3_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m3_s9_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S9_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s10_sel: begin
                              m3_nxt_st[48:0] = m3_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m3_latch_cmd = m3_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m3_s10_cmd_cur = m3_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m3_s10_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S10_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s11_sel: begin
                              m3_nxt_st[48:0] = m3_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m3_latch_cmd = m3_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m3_s11_cmd_cur = m3_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m3_s11_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S11_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             default: begin
                             m3_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m3_nxt_st[48:0] = S_S1_DATA;
end
  S_S2_CMD: begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = s2_hready ? 1'b1 : 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       m3_nxt_st[48:0] = s2_hready  ? S_S2_DATA : S_S2_CMD;
  end
  S_S2_DATA:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b1;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       if(s2_hready)
         begin
           case(1'b1)
             m3_s0_sel: begin
                              m3_nxt_st[48:0] = m3_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m3_latch_cmd = m3_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m3_s0_cmd_cur = m3_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m3_s0_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S0_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s1_sel: begin
                              m3_nxt_st[48:0] = m3_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m3_latch_cmd = m3_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m3_s1_cmd_cur = m3_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m3_s1_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S1_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s2_sel: begin
                              m3_nxt_st[48:0] = S_S2_DATA;
                              m3_s2_cmd_cur = 1'b1;
                             end
             m3_s2_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S2_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s3_sel: begin
                              m3_nxt_st[48:0] = m3_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m3_latch_cmd = m3_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m3_s3_cmd_cur = m3_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m3_s3_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S3_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s4_sel: begin
                              m3_nxt_st[48:0] = m3_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m3_latch_cmd = m3_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m3_s4_cmd_cur = m3_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m3_s4_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S4_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s5_sel: begin
                              m3_nxt_st[48:0] = m3_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m3_latch_cmd = m3_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m3_s5_cmd_cur = m3_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m3_s5_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S5_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s6_sel: begin
                              m3_nxt_st[48:0] = m3_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m3_latch_cmd = m3_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m3_s6_cmd_cur = m3_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m3_s6_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S6_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s7_sel: begin
                              m3_nxt_st[48:0] = m3_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m3_latch_cmd = m3_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m3_s7_cmd_cur = m3_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m3_s7_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S7_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s8_sel: begin
                              m3_nxt_st[48:0] = m3_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m3_latch_cmd = m3_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m3_s8_cmd_cur = m3_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m3_s8_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S8_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s9_sel: begin
                              m3_nxt_st[48:0] = m3_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m3_latch_cmd = m3_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m3_s9_cmd_cur = m3_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m3_s9_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S9_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s10_sel: begin
                              m3_nxt_st[48:0] = m3_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m3_latch_cmd = m3_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m3_s10_cmd_cur = m3_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m3_s10_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S10_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s11_sel: begin
                              m3_nxt_st[48:0] = m3_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m3_latch_cmd = m3_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m3_s11_cmd_cur = m3_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m3_s11_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S11_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             default: begin
                             m3_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m3_nxt_st[48:0] = S_S2_DATA;
end
  S_S3_CMD: begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = s3_hready ? 1'b1 : 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       m3_nxt_st[48:0] = s3_hready  ? S_S3_DATA : S_S3_CMD;
  end
  S_S3_DATA:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b1;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       if(s3_hready)
         begin
           case(1'b1)
             m3_s0_sel: begin
                              m3_nxt_st[48:0] = m3_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m3_latch_cmd = m3_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m3_s0_cmd_cur = m3_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m3_s0_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S0_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s1_sel: begin
                              m3_nxt_st[48:0] = m3_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m3_latch_cmd = m3_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m3_s1_cmd_cur = m3_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m3_s1_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S1_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s2_sel: begin
                              m3_nxt_st[48:0] = m3_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m3_latch_cmd = m3_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m3_s2_cmd_cur = m3_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m3_s2_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S2_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s3_sel: begin
                              m3_nxt_st[48:0] = S_S3_DATA;
                              m3_s3_cmd_cur = 1'b1;
                             end
             m3_s3_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S3_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s4_sel: begin
                              m3_nxt_st[48:0] = m3_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m3_latch_cmd = m3_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m3_s4_cmd_cur = m3_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m3_s4_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S4_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s5_sel: begin
                              m3_nxt_st[48:0] = m3_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m3_latch_cmd = m3_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m3_s5_cmd_cur = m3_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m3_s5_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S5_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s6_sel: begin
                              m3_nxt_st[48:0] = m3_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m3_latch_cmd = m3_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m3_s6_cmd_cur = m3_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m3_s6_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S6_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s7_sel: begin
                              m3_nxt_st[48:0] = m3_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m3_latch_cmd = m3_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m3_s7_cmd_cur = m3_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m3_s7_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S7_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s8_sel: begin
                              m3_nxt_st[48:0] = m3_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m3_latch_cmd = m3_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m3_s8_cmd_cur = m3_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m3_s8_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S8_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s9_sel: begin
                              m3_nxt_st[48:0] = m3_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m3_latch_cmd = m3_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m3_s9_cmd_cur = m3_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m3_s9_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S9_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s10_sel: begin
                              m3_nxt_st[48:0] = m3_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m3_latch_cmd = m3_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m3_s10_cmd_cur = m3_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m3_s10_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S10_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s11_sel: begin
                              m3_nxt_st[48:0] = m3_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m3_latch_cmd = m3_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m3_s11_cmd_cur = m3_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m3_s11_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S11_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             default: begin
                             m3_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m3_nxt_st[48:0] = S_S3_DATA;
end
  S_S4_CMD: begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = s4_hready ? 1'b1 : 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       m3_nxt_st[48:0] = s4_hready  ? S_S4_DATA : S_S4_CMD;
  end
  S_S4_DATA:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b1;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       if(s4_hready)
         begin
           case(1'b1)
             m3_s0_sel: begin
                              m3_nxt_st[48:0] = m3_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m3_latch_cmd = m3_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m3_s0_cmd_cur = m3_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m3_s0_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S0_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s1_sel: begin
                              m3_nxt_st[48:0] = m3_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m3_latch_cmd = m3_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m3_s1_cmd_cur = m3_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m3_s1_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S1_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s2_sel: begin
                              m3_nxt_st[48:0] = m3_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m3_latch_cmd = m3_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m3_s2_cmd_cur = m3_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m3_s2_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S2_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s3_sel: begin
                              m3_nxt_st[48:0] = m3_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m3_latch_cmd = m3_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m3_s3_cmd_cur = m3_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m3_s3_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S3_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s4_sel: begin
                              m3_nxt_st[48:0] = S_S4_DATA;
                              m3_s4_cmd_cur = 1'b1;
                             end
             m3_s4_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S4_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s5_sel: begin
                              m3_nxt_st[48:0] = m3_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m3_latch_cmd = m3_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m3_s5_cmd_cur = m3_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m3_s5_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S5_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s6_sel: begin
                              m3_nxt_st[48:0] = m3_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m3_latch_cmd = m3_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m3_s6_cmd_cur = m3_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m3_s6_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S6_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s7_sel: begin
                              m3_nxt_st[48:0] = m3_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m3_latch_cmd = m3_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m3_s7_cmd_cur = m3_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m3_s7_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S7_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s8_sel: begin
                              m3_nxt_st[48:0] = m3_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m3_latch_cmd = m3_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m3_s8_cmd_cur = m3_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m3_s8_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S8_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s9_sel: begin
                              m3_nxt_st[48:0] = m3_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m3_latch_cmd = m3_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m3_s9_cmd_cur = m3_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m3_s9_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S9_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s10_sel: begin
                              m3_nxt_st[48:0] = m3_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m3_latch_cmd = m3_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m3_s10_cmd_cur = m3_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m3_s10_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S10_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s11_sel: begin
                              m3_nxt_st[48:0] = m3_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m3_latch_cmd = m3_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m3_s11_cmd_cur = m3_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m3_s11_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S11_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             default: begin
                             m3_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m3_nxt_st[48:0] = S_S4_DATA;
end
  S_S5_CMD: begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = s5_hready ? 1'b1 : 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       m3_nxt_st[48:0] = s5_hready  ? S_S5_DATA : S_S5_CMD;
  end
  S_S5_DATA:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b1;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       if(s5_hready)
         begin
           case(1'b1)
             m3_s0_sel: begin
                              m3_nxt_st[48:0] = m3_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m3_latch_cmd = m3_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m3_s0_cmd_cur = m3_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m3_s0_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S0_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s1_sel: begin
                              m3_nxt_st[48:0] = m3_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m3_latch_cmd = m3_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m3_s1_cmd_cur = m3_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m3_s1_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S1_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s2_sel: begin
                              m3_nxt_st[48:0] = m3_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m3_latch_cmd = m3_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m3_s2_cmd_cur = m3_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m3_s2_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S2_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s3_sel: begin
                              m3_nxt_st[48:0] = m3_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m3_latch_cmd = m3_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m3_s3_cmd_cur = m3_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m3_s3_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S3_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s4_sel: begin
                              m3_nxt_st[48:0] = m3_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m3_latch_cmd = m3_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m3_s4_cmd_cur = m3_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m3_s4_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S4_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s5_sel: begin
                              m3_nxt_st[48:0] = S_S5_DATA;
                              m3_s5_cmd_cur = 1'b1;
                             end
             m3_s5_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S5_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s6_sel: begin
                              m3_nxt_st[48:0] = m3_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m3_latch_cmd = m3_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m3_s6_cmd_cur = m3_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m3_s6_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S6_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s7_sel: begin
                              m3_nxt_st[48:0] = m3_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m3_latch_cmd = m3_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m3_s7_cmd_cur = m3_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m3_s7_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S7_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s8_sel: begin
                              m3_nxt_st[48:0] = m3_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m3_latch_cmd = m3_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m3_s8_cmd_cur = m3_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m3_s8_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S8_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s9_sel: begin
                              m3_nxt_st[48:0] = m3_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m3_latch_cmd = m3_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m3_s9_cmd_cur = m3_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m3_s9_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S9_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s10_sel: begin
                              m3_nxt_st[48:0] = m3_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m3_latch_cmd = m3_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m3_s10_cmd_cur = m3_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m3_s10_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S10_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s11_sel: begin
                              m3_nxt_st[48:0] = m3_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m3_latch_cmd = m3_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m3_s11_cmd_cur = m3_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m3_s11_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S11_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             default: begin
                             m3_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m3_nxt_st[48:0] = S_S5_DATA;
end
  S_S6_CMD: begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = s6_hready ? 1'b1 : 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       m3_nxt_st[48:0] = s6_hready  ? S_S6_DATA : S_S6_CMD;
  end
  S_S6_DATA:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b1;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       if(s6_hready)
         begin
           case(1'b1)
             m3_s0_sel: begin
                              m3_nxt_st[48:0] = m3_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m3_latch_cmd = m3_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m3_s0_cmd_cur = m3_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m3_s0_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S0_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s1_sel: begin
                              m3_nxt_st[48:0] = m3_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m3_latch_cmd = m3_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m3_s1_cmd_cur = m3_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m3_s1_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S1_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s2_sel: begin
                              m3_nxt_st[48:0] = m3_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m3_latch_cmd = m3_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m3_s2_cmd_cur = m3_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m3_s2_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S2_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s3_sel: begin
                              m3_nxt_st[48:0] = m3_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m3_latch_cmd = m3_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m3_s3_cmd_cur = m3_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m3_s3_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S3_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s4_sel: begin
                              m3_nxt_st[48:0] = m3_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m3_latch_cmd = m3_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m3_s4_cmd_cur = m3_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m3_s4_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S4_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s5_sel: begin
                              m3_nxt_st[48:0] = m3_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m3_latch_cmd = m3_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m3_s5_cmd_cur = m3_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m3_s5_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S5_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s6_sel: begin
                              m3_nxt_st[48:0] = S_S6_DATA;
                              m3_s6_cmd_cur = 1'b1;
                             end
             m3_s6_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S6_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s7_sel: begin
                              m3_nxt_st[48:0] = m3_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m3_latch_cmd = m3_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m3_s7_cmd_cur = m3_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m3_s7_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S7_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s8_sel: begin
                              m3_nxt_st[48:0] = m3_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m3_latch_cmd = m3_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m3_s8_cmd_cur = m3_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m3_s8_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S8_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s9_sel: begin
                              m3_nxt_st[48:0] = m3_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m3_latch_cmd = m3_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m3_s9_cmd_cur = m3_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m3_s9_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S9_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s10_sel: begin
                              m3_nxt_st[48:0] = m3_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m3_latch_cmd = m3_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m3_s10_cmd_cur = m3_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m3_s10_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S10_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s11_sel: begin
                              m3_nxt_st[48:0] = m3_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m3_latch_cmd = m3_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m3_s11_cmd_cur = m3_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m3_s11_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S11_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             default: begin
                             m3_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m3_nxt_st[48:0] = S_S6_DATA;
end
  S_S7_CMD: begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = s7_hready ? 1'b1 : 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       m3_nxt_st[48:0] = s7_hready  ? S_S7_DATA : S_S7_CMD;
  end
  S_S7_DATA:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b1;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       if(s7_hready)
         begin
           case(1'b1)
             m3_s0_sel: begin
                              m3_nxt_st[48:0] = m3_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m3_latch_cmd = m3_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m3_s0_cmd_cur = m3_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m3_s0_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S0_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s1_sel: begin
                              m3_nxt_st[48:0] = m3_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m3_latch_cmd = m3_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m3_s1_cmd_cur = m3_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m3_s1_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S1_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s2_sel: begin
                              m3_nxt_st[48:0] = m3_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m3_latch_cmd = m3_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m3_s2_cmd_cur = m3_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m3_s2_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S2_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s3_sel: begin
                              m3_nxt_st[48:0] = m3_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m3_latch_cmd = m3_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m3_s3_cmd_cur = m3_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m3_s3_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S3_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s4_sel: begin
                              m3_nxt_st[48:0] = m3_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m3_latch_cmd = m3_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m3_s4_cmd_cur = m3_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m3_s4_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S4_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s5_sel: begin
                              m3_nxt_st[48:0] = m3_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m3_latch_cmd = m3_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m3_s5_cmd_cur = m3_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m3_s5_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S5_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s6_sel: begin
                              m3_nxt_st[48:0] = m3_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m3_latch_cmd = m3_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m3_s6_cmd_cur = m3_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m3_s6_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S6_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s7_sel: begin
                              m3_nxt_st[48:0] = S_S7_DATA;
                              m3_s7_cmd_cur = 1'b1;
                             end
             m3_s7_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S7_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s8_sel: begin
                              m3_nxt_st[48:0] = m3_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m3_latch_cmd = m3_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m3_s8_cmd_cur = m3_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m3_s8_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S8_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s9_sel: begin
                              m3_nxt_st[48:0] = m3_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m3_latch_cmd = m3_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m3_s9_cmd_cur = m3_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m3_s9_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S9_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s10_sel: begin
                              m3_nxt_st[48:0] = m3_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m3_latch_cmd = m3_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m3_s10_cmd_cur = m3_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m3_s10_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S10_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s11_sel: begin
                              m3_nxt_st[48:0] = m3_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m3_latch_cmd = m3_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m3_s11_cmd_cur = m3_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m3_s11_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S11_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             default: begin
                             m3_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m3_nxt_st[48:0] = S_S7_DATA;
end
  S_S8_CMD: begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = s8_hready ? 1'b1 : 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       m3_nxt_st[48:0] = s8_hready  ? S_S8_DATA : S_S8_CMD;
  end
  S_S8_DATA:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b1;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       if(s8_hready)
         begin
           case(1'b1)
             m3_s0_sel: begin
                              m3_nxt_st[48:0] = m3_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m3_latch_cmd = m3_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m3_s0_cmd_cur = m3_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m3_s0_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S0_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s1_sel: begin
                              m3_nxt_st[48:0] = m3_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m3_latch_cmd = m3_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m3_s1_cmd_cur = m3_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m3_s1_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S1_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s2_sel: begin
                              m3_nxt_st[48:0] = m3_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m3_latch_cmd = m3_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m3_s2_cmd_cur = m3_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m3_s2_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S2_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s3_sel: begin
                              m3_nxt_st[48:0] = m3_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m3_latch_cmd = m3_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m3_s3_cmd_cur = m3_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m3_s3_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S3_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s4_sel: begin
                              m3_nxt_st[48:0] = m3_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m3_latch_cmd = m3_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m3_s4_cmd_cur = m3_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m3_s4_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S4_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s5_sel: begin
                              m3_nxt_st[48:0] = m3_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m3_latch_cmd = m3_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m3_s5_cmd_cur = m3_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m3_s5_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S5_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s6_sel: begin
                              m3_nxt_st[48:0] = m3_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m3_latch_cmd = m3_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m3_s6_cmd_cur = m3_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m3_s6_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S6_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s7_sel: begin
                              m3_nxt_st[48:0] = m3_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m3_latch_cmd = m3_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m3_s7_cmd_cur = m3_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m3_s7_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S7_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s8_sel: begin
                              m3_nxt_st[48:0] = S_S8_DATA;
                              m3_s8_cmd_cur = 1'b1;
                             end
             m3_s8_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S8_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s9_sel: begin
                              m3_nxt_st[48:0] = m3_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m3_latch_cmd = m3_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m3_s9_cmd_cur = m3_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m3_s9_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S9_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s10_sel: begin
                              m3_nxt_st[48:0] = m3_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m3_latch_cmd = m3_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m3_s10_cmd_cur = m3_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m3_s10_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S10_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s11_sel: begin
                              m3_nxt_st[48:0] = m3_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m3_latch_cmd = m3_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m3_s11_cmd_cur = m3_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m3_s11_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S11_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             default: begin
                             m3_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m3_nxt_st[48:0] = S_S8_DATA;
end
  S_S9_CMD: begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = s9_hready ? 1'b1 : 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       m3_nxt_st[48:0] = s9_hready  ? S_S9_DATA : S_S9_CMD;
  end
  S_S9_DATA:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b1;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       if(s9_hready)
         begin
           case(1'b1)
             m3_s0_sel: begin
                              m3_nxt_st[48:0] = m3_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m3_latch_cmd = m3_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m3_s0_cmd_cur = m3_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m3_s0_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S0_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s1_sel: begin
                              m3_nxt_st[48:0] = m3_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m3_latch_cmd = m3_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m3_s1_cmd_cur = m3_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m3_s1_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S1_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s2_sel: begin
                              m3_nxt_st[48:0] = m3_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m3_latch_cmd = m3_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m3_s2_cmd_cur = m3_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m3_s2_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S2_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s3_sel: begin
                              m3_nxt_st[48:0] = m3_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m3_latch_cmd = m3_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m3_s3_cmd_cur = m3_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m3_s3_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S3_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s4_sel: begin
                              m3_nxt_st[48:0] = m3_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m3_latch_cmd = m3_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m3_s4_cmd_cur = m3_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m3_s4_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S4_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s5_sel: begin
                              m3_nxt_st[48:0] = m3_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m3_latch_cmd = m3_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m3_s5_cmd_cur = m3_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m3_s5_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S5_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s6_sel: begin
                              m3_nxt_st[48:0] = m3_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m3_latch_cmd = m3_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m3_s6_cmd_cur = m3_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m3_s6_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S6_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s7_sel: begin
                              m3_nxt_st[48:0] = m3_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m3_latch_cmd = m3_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m3_s7_cmd_cur = m3_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m3_s7_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S7_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s8_sel: begin
                              m3_nxt_st[48:0] = m3_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m3_latch_cmd = m3_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m3_s8_cmd_cur = m3_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m3_s8_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S8_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s9_sel: begin
                              m3_nxt_st[48:0] = S_S9_DATA;
                              m3_s9_cmd_cur = 1'b1;
                             end
             m3_s9_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S9_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s10_sel: begin
                              m3_nxt_st[48:0] = m3_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m3_latch_cmd = m3_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m3_s10_cmd_cur = m3_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m3_s10_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S10_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s11_sel: begin
                              m3_nxt_st[48:0] = m3_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m3_latch_cmd = m3_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m3_s11_cmd_cur = m3_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m3_s11_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S11_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             default: begin
                             m3_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m3_nxt_st[48:0] = S_S9_DATA;
end
  S_S10_CMD: begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = s10_hready ? 1'b1 : 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       m3_nxt_st[48:0] = s10_hready  ? S_S10_DATA : S_S10_CMD;
  end
  S_S10_DATA:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b1;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       if(s10_hready)
         begin
           case(1'b1)
             m3_s0_sel: begin
                              m3_nxt_st[48:0] = m3_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m3_latch_cmd = m3_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m3_s0_cmd_cur = m3_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m3_s0_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S0_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s1_sel: begin
                              m3_nxt_st[48:0] = m3_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m3_latch_cmd = m3_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m3_s1_cmd_cur = m3_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m3_s1_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S1_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s2_sel: begin
                              m3_nxt_st[48:0] = m3_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m3_latch_cmd = m3_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m3_s2_cmd_cur = m3_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m3_s2_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S2_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s3_sel: begin
                              m3_nxt_st[48:0] = m3_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m3_latch_cmd = m3_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m3_s3_cmd_cur = m3_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m3_s3_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S3_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s4_sel: begin
                              m3_nxt_st[48:0] = m3_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m3_latch_cmd = m3_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m3_s4_cmd_cur = m3_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m3_s4_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S4_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s5_sel: begin
                              m3_nxt_st[48:0] = m3_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m3_latch_cmd = m3_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m3_s5_cmd_cur = m3_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m3_s5_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S5_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s6_sel: begin
                              m3_nxt_st[48:0] = m3_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m3_latch_cmd = m3_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m3_s6_cmd_cur = m3_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m3_s6_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S6_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s7_sel: begin
                              m3_nxt_st[48:0] = m3_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m3_latch_cmd = m3_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m3_s7_cmd_cur = m3_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m3_s7_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S7_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s8_sel: begin
                              m3_nxt_st[48:0] = m3_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m3_latch_cmd = m3_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m3_s8_cmd_cur = m3_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m3_s8_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S8_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s9_sel: begin
                              m3_nxt_st[48:0] = m3_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m3_latch_cmd = m3_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m3_s9_cmd_cur = m3_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m3_s9_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S9_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s10_sel: begin
                              m3_nxt_st[48:0] = S_S10_DATA;
                              m3_s10_cmd_cur = 1'b1;
                             end
             m3_s10_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S10_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s11_sel: begin
                              m3_nxt_st[48:0] = m3_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m3_latch_cmd = m3_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m3_s11_cmd_cur = m3_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m3_s11_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S11_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             default: begin
                             m3_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m3_nxt_st[48:0] = S_S10_DATA;
end
  S_S11_CMD: begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = s11_hready ? 1'b1 : 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b0;
       m3_nxt_st[48:0] = s11_hready  ? S_S11_DATA : S_S11_CMD;
  end
  S_S11_DATA:begin
       m3_latch_cmd = 1'b0;
       m3_s0_cmd_last = 1'b0;
       m3_s0_cmd_cur = 1'b0;
       m3_s0_data = 1'b0;
       m3_s1_cmd_last = 1'b0;
       m3_s1_cmd_cur = 1'b0;
       m3_s1_data = 1'b0;
       m3_s2_cmd_last = 1'b0;
       m3_s2_cmd_cur = 1'b0;
       m3_s2_data = 1'b0;
       m3_s3_cmd_last = 1'b0;
       m3_s3_cmd_cur = 1'b0;
       m3_s3_data = 1'b0;
       m3_s4_cmd_last = 1'b0;
       m3_s4_cmd_cur = 1'b0;
       m3_s4_data = 1'b0;
       m3_s5_cmd_last = 1'b0;
       m3_s5_cmd_cur = 1'b0;
       m3_s5_data = 1'b0;
       m3_s6_cmd_last = 1'b0;
       m3_s6_cmd_cur = 1'b0;
       m3_s6_data = 1'b0;
       m3_s7_cmd_last = 1'b0;
       m3_s7_cmd_cur = 1'b0;
       m3_s7_data = 1'b0;
       m3_s8_cmd_last = 1'b0;
       m3_s8_cmd_cur = 1'b0;
       m3_s8_data = 1'b0;
       m3_s9_cmd_last = 1'b0;
       m3_s9_cmd_cur = 1'b0;
       m3_s9_data = 1'b0;
       m3_s10_cmd_last = 1'b0;
       m3_s10_cmd_cur = 1'b0;
       m3_s10_data = 1'b0;
       m3_s11_cmd_last = 1'b0;
       m3_s11_cmd_cur = 1'b0;
       m3_s11_data = 1'b1;
       if(s11_hready)
         begin
           case(1'b1)
             m3_s0_sel: begin
                              m3_nxt_st[48:0] = m3_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m3_latch_cmd = m3_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m3_s0_cmd_cur = m3_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m3_s0_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S0_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s1_sel: begin
                              m3_nxt_st[48:0] = m3_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m3_latch_cmd = m3_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m3_s1_cmd_cur = m3_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m3_s1_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S1_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s2_sel: begin
                              m3_nxt_st[48:0] = m3_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m3_latch_cmd = m3_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m3_s2_cmd_cur = m3_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m3_s2_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S2_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s3_sel: begin
                              m3_nxt_st[48:0] = m3_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m3_latch_cmd = m3_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m3_s3_cmd_cur = m3_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m3_s3_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S3_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s4_sel: begin
                              m3_nxt_st[48:0] = m3_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m3_latch_cmd = m3_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m3_s4_cmd_cur = m3_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m3_s4_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S4_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s5_sel: begin
                              m3_nxt_st[48:0] = m3_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m3_latch_cmd = m3_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m3_s5_cmd_cur = m3_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m3_s5_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S5_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s6_sel: begin
                              m3_nxt_st[48:0] = m3_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m3_latch_cmd = m3_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m3_s6_cmd_cur = m3_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m3_s6_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S6_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s7_sel: begin
                              m3_nxt_st[48:0] = m3_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m3_latch_cmd = m3_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m3_s7_cmd_cur = m3_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m3_s7_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S7_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s8_sel: begin
                              m3_nxt_st[48:0] = m3_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m3_latch_cmd = m3_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m3_s8_cmd_cur = m3_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m3_s8_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S8_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s9_sel: begin
                              m3_nxt_st[48:0] = m3_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m3_latch_cmd = m3_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m3_s9_cmd_cur = m3_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m3_s9_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S9_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s10_sel: begin
                              m3_nxt_st[48:0] = m3_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m3_latch_cmd = m3_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m3_s10_cmd_cur = m3_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m3_s10_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S10_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             m3_s11_sel: begin
                              m3_nxt_st[48:0] = S_S11_DATA;
                              m3_s11_cmd_cur = 1'b1;
                             end
             m3_s11_wt_sel: begin
                                 m3_nxt_st[48:0] = S_S11_GNT;
                                 m3_latch_cmd = 1'b1;
                               end
             default: begin
                             m3_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m3_nxt_st[48:0] = S_S11_DATA;
end
  default: begin
             m3_latch_cmd = 1'b0;
             m3_s0_cmd_last = 1'b0;
             m3_s0_cmd_cur = 1'b0;
             m3_s0_data = 1'b0;
             m3_s1_cmd_last = 1'b0;
             m3_s1_cmd_cur = 1'b0;
             m3_s1_data = 1'b0;
             m3_s2_cmd_last = 1'b0;
             m3_s2_cmd_cur = 1'b0;
             m3_s2_data = 1'b0;
             m3_s3_cmd_last = 1'b0;
             m3_s3_cmd_cur = 1'b0;
             m3_s3_data = 1'b0;
             m3_s4_cmd_last = 1'b0;
             m3_s4_cmd_cur = 1'b0;
             m3_s4_data = 1'b0;
             m3_s5_cmd_last = 1'b0;
             m3_s5_cmd_cur = 1'b0;
             m3_s5_data = 1'b0;
             m3_s6_cmd_last = 1'b0;
             m3_s6_cmd_cur = 1'b0;
             m3_s6_data = 1'b0;
             m3_s7_cmd_last = 1'b0;
             m3_s7_cmd_cur = 1'b0;
             m3_s7_data = 1'b0;
             m3_s8_cmd_last = 1'b0;
             m3_s8_cmd_cur = 1'b0;
             m3_s8_data = 1'b0;
             m3_s9_cmd_last = 1'b0;
             m3_s9_cmd_cur = 1'b0;
             m3_s9_data = 1'b0;
             m3_s10_cmd_last = 1'b0;
             m3_s10_cmd_cur = 1'b0;
             m3_s10_data = 1'b0;
             m3_s11_cmd_last = 1'b0;
             m3_s11_cmd_cur = 1'b0;
             m3_s11_data = 1'b0;
             m3_nxt_st[48:0] = S_IDLE;
  end
endcase
end
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
       m4_cur_st[48:0] <= S_IDLE;
    else
       m4_cur_st[48:0] <= m4_nxt_st[48:0];
  end
always @ (*)
begin
case(m4_cur_st[48:0])
  S_IDLE:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       case(1'b1)
         m4_s0_sel: begin
                          m4_nxt_st[48:0] = m4_s0_hld ? S_S0_WAIT : (s0_hready ? S_S0_DATA : S_S0_CMD);
                          m4_latch_cmd = m4_s0_hld ? 1'b1 : (s0_hready ? 1'b0 : 1'b1);
                          m4_s0_cmd_cur = m4_s0_hld ? 1'b0 : (s0_hready ? 1'b1 : 1'b0);
                        end
         m4_s0_wt_sel: begin
                             m4_nxt_st[48:0] = S_S0_GNT;
                             m4_latch_cmd = 1'b1;
                           end
         m4_s1_sel: begin
                          m4_nxt_st[48:0] = m4_s1_hld ? S_S1_WAIT : (s1_hready ? S_S1_DATA : S_S1_CMD);
                          m4_latch_cmd = m4_s1_hld ? 1'b1 : (s1_hready ? 1'b0 : 1'b1);
                          m4_s1_cmd_cur = m4_s1_hld ? 1'b0 : (s1_hready ? 1'b1 : 1'b0);
                        end
         m4_s1_wt_sel: begin
                             m4_nxt_st[48:0] = S_S1_GNT;
                             m4_latch_cmd = 1'b1;
                           end
         m4_s2_sel: begin
                          m4_nxt_st[48:0] = m4_s2_hld ? S_S2_WAIT : (s2_hready ? S_S2_DATA : S_S2_CMD);
                          m4_latch_cmd = m4_s2_hld ? 1'b1 : (s2_hready ? 1'b0 : 1'b1);
                          m4_s2_cmd_cur = m4_s2_hld ? 1'b0 : (s2_hready ? 1'b1 : 1'b0);
                        end
         m4_s2_wt_sel: begin
                             m4_nxt_st[48:0] = S_S2_GNT;
                             m4_latch_cmd = 1'b1;
                           end
         m4_s3_sel: begin
                          m4_nxt_st[48:0] = m4_s3_hld ? S_S3_WAIT : (s3_hready ? S_S3_DATA : S_S3_CMD);
                          m4_latch_cmd = m4_s3_hld ? 1'b1 : (s3_hready ? 1'b0 : 1'b1);
                          m4_s3_cmd_cur = m4_s3_hld ? 1'b0 : (s3_hready ? 1'b1 : 1'b0);
                        end
         m4_s3_wt_sel: begin
                             m4_nxt_st[48:0] = S_S3_GNT;
                             m4_latch_cmd = 1'b1;
                           end
         m4_s4_sel: begin
                          m4_nxt_st[48:0] = m4_s4_hld ? S_S4_WAIT : (s4_hready ? S_S4_DATA : S_S4_CMD);
                          m4_latch_cmd = m4_s4_hld ? 1'b1 : (s4_hready ? 1'b0 : 1'b1);
                          m4_s4_cmd_cur = m4_s4_hld ? 1'b0 : (s4_hready ? 1'b1 : 1'b0);
                        end
         m4_s4_wt_sel: begin
                             m4_nxt_st[48:0] = S_S4_GNT;
                             m4_latch_cmd = 1'b1;
                           end
         m4_s5_sel: begin
                          m4_nxt_st[48:0] = m4_s5_hld ? S_S5_WAIT : (s5_hready ? S_S5_DATA : S_S5_CMD);
                          m4_latch_cmd = m4_s5_hld ? 1'b1 : (s5_hready ? 1'b0 : 1'b1);
                          m4_s5_cmd_cur = m4_s5_hld ? 1'b0 : (s5_hready ? 1'b1 : 1'b0);
                        end
         m4_s5_wt_sel: begin
                             m4_nxt_st[48:0] = S_S5_GNT;
                             m4_latch_cmd = 1'b1;
                           end
         m4_s6_sel: begin
                          m4_nxt_st[48:0] = m4_s6_hld ? S_S6_WAIT : (s6_hready ? S_S6_DATA : S_S6_CMD);
                          m4_latch_cmd = m4_s6_hld ? 1'b1 : (s6_hready ? 1'b0 : 1'b1);
                          m4_s6_cmd_cur = m4_s6_hld ? 1'b0 : (s6_hready ? 1'b1 : 1'b0);
                        end
         m4_s6_wt_sel: begin
                             m4_nxt_st[48:0] = S_S6_GNT;
                             m4_latch_cmd = 1'b1;
                           end
         m4_s7_sel: begin
                          m4_nxt_st[48:0] = m4_s7_hld ? S_S7_WAIT : (s7_hready ? S_S7_DATA : S_S7_CMD);
                          m4_latch_cmd = m4_s7_hld ? 1'b1 : (s7_hready ? 1'b0 : 1'b1);
                          m4_s7_cmd_cur = m4_s7_hld ? 1'b0 : (s7_hready ? 1'b1 : 1'b0);
                        end
         m4_s7_wt_sel: begin
                             m4_nxt_st[48:0] = S_S7_GNT;
                             m4_latch_cmd = 1'b1;
                           end
         m4_s8_sel: begin
                          m4_nxt_st[48:0] = m4_s8_hld ? S_S8_WAIT : (s8_hready ? S_S8_DATA : S_S8_CMD);
                          m4_latch_cmd = m4_s8_hld ? 1'b1 : (s8_hready ? 1'b0 : 1'b1);
                          m4_s8_cmd_cur = m4_s8_hld ? 1'b0 : (s8_hready ? 1'b1 : 1'b0);
                        end
         m4_s8_wt_sel: begin
                             m4_nxt_st[48:0] = S_S8_GNT;
                             m4_latch_cmd = 1'b1;
                           end
         m4_s9_sel: begin
                          m4_nxt_st[48:0] = m4_s9_hld ? S_S9_WAIT : (s9_hready ? S_S9_DATA : S_S9_CMD);
                          m4_latch_cmd = m4_s9_hld ? 1'b1 : (s9_hready ? 1'b0 : 1'b1);
                          m4_s9_cmd_cur = m4_s9_hld ? 1'b0 : (s9_hready ? 1'b1 : 1'b0);
                        end
         m4_s9_wt_sel: begin
                             m4_nxt_st[48:0] = S_S9_GNT;
                             m4_latch_cmd = 1'b1;
                           end
         m4_s10_sel: begin
                          m4_nxt_st[48:0] = m4_s10_hld ? S_S10_WAIT : (s10_hready ? S_S10_DATA : S_S10_CMD);
                          m4_latch_cmd = m4_s10_hld ? 1'b1 : (s10_hready ? 1'b0 : 1'b1);
                          m4_s10_cmd_cur = m4_s10_hld ? 1'b0 : (s10_hready ? 1'b1 : 1'b0);
                        end
         m4_s10_wt_sel: begin
                             m4_nxt_st[48:0] = S_S10_GNT;
                             m4_latch_cmd = 1'b1;
                           end
         m4_s11_sel: begin
                          m4_nxt_st[48:0] = m4_s11_hld ? S_S11_WAIT : (s11_hready ? S_S11_DATA : S_S11_CMD);
                          m4_latch_cmd = m4_s11_hld ? 1'b1 : (s11_hready ? 1'b0 : 1'b1);
                          m4_s11_cmd_cur = m4_s11_hld ? 1'b0 : (s11_hready ? 1'b1 : 1'b0);
                        end
         m4_s11_wt_sel: begin
                             m4_nxt_st[48:0] = S_S11_GNT;
                             m4_latch_cmd = 1'b1;
                           end
         default: begin
                          m4_nxt_st[48:0] = S_IDLE;
                  end
       endcase
  end
  S_S0_GNT:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       case(1'b1)
         m4_s0_sel: begin
                          m4_nxt_st[48:0] = m4_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                          m4_s0_cmd_last = m4_s0_hld ? 1'b0 : (s0_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m4_nxt_st[48:0] = S_S0_GNT;
                  end
       endcase
  end
  S_S1_GNT:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       case(1'b1)
         m4_s1_sel: begin
                          m4_nxt_st[48:0] = m4_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                          m4_s1_cmd_last = m4_s1_hld ? 1'b0 : (s1_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m4_nxt_st[48:0] = S_S1_GNT;
                  end
       endcase
  end
  S_S2_GNT:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       case(1'b1)
         m4_s2_sel: begin
                          m4_nxt_st[48:0] = m4_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                          m4_s2_cmd_last = m4_s2_hld ? 1'b0 : (s2_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m4_nxt_st[48:0] = S_S2_GNT;
                  end
       endcase
  end
  S_S3_GNT:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       case(1'b1)
         m4_s3_sel: begin
                          m4_nxt_st[48:0] = m4_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                          m4_s3_cmd_last = m4_s3_hld ? 1'b0 : (s3_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m4_nxt_st[48:0] = S_S3_GNT;
                  end
       endcase
  end
  S_S4_GNT:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       case(1'b1)
         m4_s4_sel: begin
                          m4_nxt_st[48:0] = m4_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                          m4_s4_cmd_last = m4_s4_hld ? 1'b0 : (s4_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m4_nxt_st[48:0] = S_S4_GNT;
                  end
       endcase
  end
  S_S5_GNT:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       case(1'b1)
         m4_s5_sel: begin
                          m4_nxt_st[48:0] = m4_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                          m4_s5_cmd_last = m4_s5_hld ? 1'b0 : (s5_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m4_nxt_st[48:0] = S_S5_GNT;
                  end
       endcase
  end
  S_S6_GNT:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       case(1'b1)
         m4_s6_sel: begin
                          m4_nxt_st[48:0] = m4_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                          m4_s6_cmd_last = m4_s6_hld ? 1'b0 : (s6_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m4_nxt_st[48:0] = S_S6_GNT;
                  end
       endcase
  end
  S_S7_GNT:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       case(1'b1)
         m4_s7_sel: begin
                          m4_nxt_st[48:0] = m4_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                          m4_s7_cmd_last = m4_s7_hld ? 1'b0 : (s7_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m4_nxt_st[48:0] = S_S7_GNT;
                  end
       endcase
  end
  S_S8_GNT:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       case(1'b1)
         m4_s8_sel: begin
                          m4_nxt_st[48:0] = m4_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                          m4_s8_cmd_last = m4_s8_hld ? 1'b0 : (s8_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m4_nxt_st[48:0] = S_S8_GNT;
                  end
       endcase
  end
  S_S9_GNT:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       case(1'b1)
         m4_s9_sel: begin
                          m4_nxt_st[48:0] = m4_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                          m4_s9_cmd_last = m4_s9_hld ? 1'b0 : (s9_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m4_nxt_st[48:0] = S_S9_GNT;
                  end
       endcase
  end
  S_S10_GNT:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       case(1'b1)
         m4_s10_sel: begin
                          m4_nxt_st[48:0] = m4_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                          m4_s10_cmd_last = m4_s10_hld ? 1'b0 : (s10_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m4_nxt_st[48:0] = S_S10_GNT;
                  end
       endcase
  end
  S_S11_GNT:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       case(1'b1)
         m4_s11_sel: begin
                          m4_nxt_st[48:0] = m4_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                          m4_s11_cmd_last = m4_s11_hld ? 1'b0 : (s11_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m4_nxt_st[48:0] = S_S11_GNT;
                  end
       endcase
  end
  S_S0_WAIT:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       case(1'b1)
         ~m4_s0_hld: begin
                          m4_nxt_st[48:0] = m4_s0_wt_sel ? S_S0_GNT : s0_hready ? S_S0_DATA : S_S0_CMD;
                          m4_s0_cmd_last = m4_s0_wt_sel ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m4_nxt_st[48:0] = S_S0_WAIT;
                  end
       endcase
  end
  S_S1_WAIT:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       case(1'b1)
         ~m4_s1_hld: begin
                          m4_nxt_st[48:0] = m4_s1_wt_sel ? S_S1_GNT : s1_hready ? S_S1_DATA : S_S1_CMD;
                          m4_s1_cmd_last = m4_s1_wt_sel ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m4_nxt_st[48:0] = S_S1_WAIT;
                  end
       endcase
  end
  S_S2_WAIT:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       case(1'b1)
         ~m4_s2_hld: begin
                          m4_nxt_st[48:0] = m4_s2_wt_sel ? S_S2_GNT : s2_hready ? S_S2_DATA : S_S2_CMD;
                          m4_s2_cmd_last = m4_s2_wt_sel ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m4_nxt_st[48:0] = S_S2_WAIT;
                  end
       endcase
  end
  S_S3_WAIT:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       case(1'b1)
         ~m4_s3_hld: begin
                          m4_nxt_st[48:0] = m4_s3_wt_sel ? S_S3_GNT : s3_hready ? S_S3_DATA : S_S3_CMD;
                          m4_s3_cmd_last = m4_s3_wt_sel ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m4_nxt_st[48:0] = S_S3_WAIT;
                  end
       endcase
  end
  S_S4_WAIT:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       case(1'b1)
         ~m4_s4_hld: begin
                          m4_nxt_st[48:0] = m4_s4_wt_sel ? S_S4_GNT : s4_hready ? S_S4_DATA : S_S4_CMD;
                          m4_s4_cmd_last = m4_s4_wt_sel ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m4_nxt_st[48:0] = S_S4_WAIT;
                  end
       endcase
  end
  S_S5_WAIT:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       case(1'b1)
         ~m4_s5_hld: begin
                          m4_nxt_st[48:0] = m4_s5_wt_sel ? S_S5_GNT : s5_hready ? S_S5_DATA : S_S5_CMD;
                          m4_s5_cmd_last = m4_s5_wt_sel ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m4_nxt_st[48:0] = S_S5_WAIT;
                  end
       endcase
  end
  S_S6_WAIT:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       case(1'b1)
         ~m4_s6_hld: begin
                          m4_nxt_st[48:0] = m4_s6_wt_sel ? S_S6_GNT : s6_hready ? S_S6_DATA : S_S6_CMD;
                          m4_s6_cmd_last = m4_s6_wt_sel ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m4_nxt_st[48:0] = S_S6_WAIT;
                  end
       endcase
  end
  S_S7_WAIT:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       case(1'b1)
         ~m4_s7_hld: begin
                          m4_nxt_st[48:0] = m4_s7_wt_sel ? S_S7_GNT : s7_hready ? S_S7_DATA : S_S7_CMD;
                          m4_s7_cmd_last = m4_s7_wt_sel ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m4_nxt_st[48:0] = S_S7_WAIT;
                  end
       endcase
  end
  S_S8_WAIT:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       case(1'b1)
         ~m4_s8_hld: begin
                          m4_nxt_st[48:0] = m4_s8_wt_sel ? S_S8_GNT : s8_hready ? S_S8_DATA : S_S8_CMD;
                          m4_s8_cmd_last = m4_s8_wt_sel ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m4_nxt_st[48:0] = S_S8_WAIT;
                  end
       endcase
  end
  S_S9_WAIT:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       case(1'b1)
         ~m4_s9_hld: begin
                          m4_nxt_st[48:0] = m4_s9_wt_sel ? S_S9_GNT : s9_hready ? S_S9_DATA : S_S9_CMD;
                          m4_s9_cmd_last = m4_s9_wt_sel ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m4_nxt_st[48:0] = S_S9_WAIT;
                  end
       endcase
  end
  S_S10_WAIT:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       case(1'b1)
         ~m4_s10_hld: begin
                          m4_nxt_st[48:0] = m4_s10_wt_sel ? S_S10_GNT : s10_hready ? S_S10_DATA : S_S10_CMD;
                          m4_s10_cmd_last = m4_s10_wt_sel ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m4_nxt_st[48:0] = S_S10_WAIT;
                  end
       endcase
  end
  S_S11_WAIT:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       case(1'b1)
         ~m4_s11_hld: begin
                          m4_nxt_st[48:0] = m4_s11_wt_sel ? S_S11_GNT : s11_hready ? S_S11_DATA : S_S11_CMD;
                          m4_s11_cmd_last = m4_s11_wt_sel ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m4_nxt_st[48:0] = S_S11_WAIT;
                  end
       endcase
  end
  S_S0_CMD: begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = s0_hready ? 1'b1 : 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       m4_nxt_st[48:0] = s0_hready  ? S_S0_DATA : S_S0_CMD;
  end
  S_S0_DATA:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b1;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       if(s0_hready)
         begin
           case(1'b1)
             m4_s0_sel: begin
                              m4_nxt_st[48:0] = S_S0_DATA;
                              m4_s0_cmd_cur = 1'b1;
                             end
             m4_s0_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S0_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s1_sel: begin
                              m4_nxt_st[48:0] = m4_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m4_latch_cmd = m4_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m4_s1_cmd_cur = m4_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m4_s1_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S1_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s2_sel: begin
                              m4_nxt_st[48:0] = m4_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m4_latch_cmd = m4_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m4_s2_cmd_cur = m4_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m4_s2_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S2_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s3_sel: begin
                              m4_nxt_st[48:0] = m4_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m4_latch_cmd = m4_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m4_s3_cmd_cur = m4_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m4_s3_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S3_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s4_sel: begin
                              m4_nxt_st[48:0] = m4_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m4_latch_cmd = m4_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m4_s4_cmd_cur = m4_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m4_s4_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S4_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s5_sel: begin
                              m4_nxt_st[48:0] = m4_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m4_latch_cmd = m4_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m4_s5_cmd_cur = m4_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m4_s5_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S5_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s6_sel: begin
                              m4_nxt_st[48:0] = m4_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m4_latch_cmd = m4_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m4_s6_cmd_cur = m4_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m4_s6_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S6_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s7_sel: begin
                              m4_nxt_st[48:0] = m4_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m4_latch_cmd = m4_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m4_s7_cmd_cur = m4_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m4_s7_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S7_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s8_sel: begin
                              m4_nxt_st[48:0] = m4_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m4_latch_cmd = m4_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m4_s8_cmd_cur = m4_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m4_s8_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S8_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s9_sel: begin
                              m4_nxt_st[48:0] = m4_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m4_latch_cmd = m4_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m4_s9_cmd_cur = m4_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m4_s9_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S9_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s10_sel: begin
                              m4_nxt_st[48:0] = m4_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m4_latch_cmd = m4_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m4_s10_cmd_cur = m4_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m4_s10_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S10_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s11_sel: begin
                              m4_nxt_st[48:0] = m4_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m4_latch_cmd = m4_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m4_s11_cmd_cur = m4_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m4_s11_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S11_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             default: begin
                             m4_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m4_nxt_st[48:0] = S_S0_DATA;
end
  S_S1_CMD: begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = s1_hready ? 1'b1 : 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       m4_nxt_st[48:0] = s1_hready  ? S_S1_DATA : S_S1_CMD;
  end
  S_S1_DATA:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b1;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       if(s1_hready)
         begin
           case(1'b1)
             m4_s0_sel: begin
                              m4_nxt_st[48:0] = m4_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m4_latch_cmd = m4_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m4_s0_cmd_cur = m4_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m4_s0_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S0_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s1_sel: begin
                              m4_nxt_st[48:0] = S_S1_DATA;
                              m4_s1_cmd_cur = 1'b1;
                             end
             m4_s1_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S1_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s2_sel: begin
                              m4_nxt_st[48:0] = m4_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m4_latch_cmd = m4_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m4_s2_cmd_cur = m4_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m4_s2_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S2_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s3_sel: begin
                              m4_nxt_st[48:0] = m4_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m4_latch_cmd = m4_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m4_s3_cmd_cur = m4_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m4_s3_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S3_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s4_sel: begin
                              m4_nxt_st[48:0] = m4_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m4_latch_cmd = m4_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m4_s4_cmd_cur = m4_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m4_s4_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S4_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s5_sel: begin
                              m4_nxt_st[48:0] = m4_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m4_latch_cmd = m4_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m4_s5_cmd_cur = m4_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m4_s5_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S5_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s6_sel: begin
                              m4_nxt_st[48:0] = m4_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m4_latch_cmd = m4_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m4_s6_cmd_cur = m4_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m4_s6_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S6_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s7_sel: begin
                              m4_nxt_st[48:0] = m4_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m4_latch_cmd = m4_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m4_s7_cmd_cur = m4_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m4_s7_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S7_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s8_sel: begin
                              m4_nxt_st[48:0] = m4_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m4_latch_cmd = m4_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m4_s8_cmd_cur = m4_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m4_s8_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S8_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s9_sel: begin
                              m4_nxt_st[48:0] = m4_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m4_latch_cmd = m4_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m4_s9_cmd_cur = m4_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m4_s9_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S9_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s10_sel: begin
                              m4_nxt_st[48:0] = m4_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m4_latch_cmd = m4_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m4_s10_cmd_cur = m4_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m4_s10_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S10_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s11_sel: begin
                              m4_nxt_st[48:0] = m4_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m4_latch_cmd = m4_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m4_s11_cmd_cur = m4_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m4_s11_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S11_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             default: begin
                             m4_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m4_nxt_st[48:0] = S_S1_DATA;
end
  S_S2_CMD: begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = s2_hready ? 1'b1 : 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       m4_nxt_st[48:0] = s2_hready  ? S_S2_DATA : S_S2_CMD;
  end
  S_S2_DATA:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b1;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       if(s2_hready)
         begin
           case(1'b1)
             m4_s0_sel: begin
                              m4_nxt_st[48:0] = m4_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m4_latch_cmd = m4_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m4_s0_cmd_cur = m4_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m4_s0_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S0_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s1_sel: begin
                              m4_nxt_st[48:0] = m4_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m4_latch_cmd = m4_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m4_s1_cmd_cur = m4_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m4_s1_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S1_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s2_sel: begin
                              m4_nxt_st[48:0] = S_S2_DATA;
                              m4_s2_cmd_cur = 1'b1;
                             end
             m4_s2_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S2_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s3_sel: begin
                              m4_nxt_st[48:0] = m4_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m4_latch_cmd = m4_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m4_s3_cmd_cur = m4_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m4_s3_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S3_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s4_sel: begin
                              m4_nxt_st[48:0] = m4_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m4_latch_cmd = m4_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m4_s4_cmd_cur = m4_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m4_s4_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S4_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s5_sel: begin
                              m4_nxt_st[48:0] = m4_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m4_latch_cmd = m4_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m4_s5_cmd_cur = m4_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m4_s5_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S5_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s6_sel: begin
                              m4_nxt_st[48:0] = m4_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m4_latch_cmd = m4_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m4_s6_cmd_cur = m4_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m4_s6_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S6_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s7_sel: begin
                              m4_nxt_st[48:0] = m4_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m4_latch_cmd = m4_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m4_s7_cmd_cur = m4_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m4_s7_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S7_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s8_sel: begin
                              m4_nxt_st[48:0] = m4_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m4_latch_cmd = m4_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m4_s8_cmd_cur = m4_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m4_s8_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S8_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s9_sel: begin
                              m4_nxt_st[48:0] = m4_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m4_latch_cmd = m4_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m4_s9_cmd_cur = m4_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m4_s9_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S9_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s10_sel: begin
                              m4_nxt_st[48:0] = m4_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m4_latch_cmd = m4_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m4_s10_cmd_cur = m4_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m4_s10_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S10_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s11_sel: begin
                              m4_nxt_st[48:0] = m4_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m4_latch_cmd = m4_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m4_s11_cmd_cur = m4_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m4_s11_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S11_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             default: begin
                             m4_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m4_nxt_st[48:0] = S_S2_DATA;
end
  S_S3_CMD: begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = s3_hready ? 1'b1 : 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       m4_nxt_st[48:0] = s3_hready  ? S_S3_DATA : S_S3_CMD;
  end
  S_S3_DATA:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b1;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       if(s3_hready)
         begin
           case(1'b1)
             m4_s0_sel: begin
                              m4_nxt_st[48:0] = m4_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m4_latch_cmd = m4_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m4_s0_cmd_cur = m4_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m4_s0_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S0_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s1_sel: begin
                              m4_nxt_st[48:0] = m4_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m4_latch_cmd = m4_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m4_s1_cmd_cur = m4_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m4_s1_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S1_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s2_sel: begin
                              m4_nxt_st[48:0] = m4_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m4_latch_cmd = m4_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m4_s2_cmd_cur = m4_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m4_s2_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S2_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s3_sel: begin
                              m4_nxt_st[48:0] = S_S3_DATA;
                              m4_s3_cmd_cur = 1'b1;
                             end
             m4_s3_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S3_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s4_sel: begin
                              m4_nxt_st[48:0] = m4_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m4_latch_cmd = m4_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m4_s4_cmd_cur = m4_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m4_s4_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S4_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s5_sel: begin
                              m4_nxt_st[48:0] = m4_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m4_latch_cmd = m4_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m4_s5_cmd_cur = m4_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m4_s5_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S5_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s6_sel: begin
                              m4_nxt_st[48:0] = m4_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m4_latch_cmd = m4_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m4_s6_cmd_cur = m4_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m4_s6_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S6_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s7_sel: begin
                              m4_nxt_st[48:0] = m4_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m4_latch_cmd = m4_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m4_s7_cmd_cur = m4_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m4_s7_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S7_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s8_sel: begin
                              m4_nxt_st[48:0] = m4_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m4_latch_cmd = m4_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m4_s8_cmd_cur = m4_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m4_s8_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S8_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s9_sel: begin
                              m4_nxt_st[48:0] = m4_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m4_latch_cmd = m4_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m4_s9_cmd_cur = m4_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m4_s9_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S9_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s10_sel: begin
                              m4_nxt_st[48:0] = m4_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m4_latch_cmd = m4_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m4_s10_cmd_cur = m4_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m4_s10_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S10_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s11_sel: begin
                              m4_nxt_st[48:0] = m4_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m4_latch_cmd = m4_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m4_s11_cmd_cur = m4_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m4_s11_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S11_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             default: begin
                             m4_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m4_nxt_st[48:0] = S_S3_DATA;
end
  S_S4_CMD: begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = s4_hready ? 1'b1 : 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       m4_nxt_st[48:0] = s4_hready  ? S_S4_DATA : S_S4_CMD;
  end
  S_S4_DATA:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b1;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       if(s4_hready)
         begin
           case(1'b1)
             m4_s0_sel: begin
                              m4_nxt_st[48:0] = m4_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m4_latch_cmd = m4_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m4_s0_cmd_cur = m4_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m4_s0_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S0_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s1_sel: begin
                              m4_nxt_st[48:0] = m4_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m4_latch_cmd = m4_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m4_s1_cmd_cur = m4_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m4_s1_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S1_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s2_sel: begin
                              m4_nxt_st[48:0] = m4_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m4_latch_cmd = m4_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m4_s2_cmd_cur = m4_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m4_s2_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S2_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s3_sel: begin
                              m4_nxt_st[48:0] = m4_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m4_latch_cmd = m4_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m4_s3_cmd_cur = m4_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m4_s3_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S3_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s4_sel: begin
                              m4_nxt_st[48:0] = S_S4_DATA;
                              m4_s4_cmd_cur = 1'b1;
                             end
             m4_s4_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S4_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s5_sel: begin
                              m4_nxt_st[48:0] = m4_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m4_latch_cmd = m4_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m4_s5_cmd_cur = m4_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m4_s5_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S5_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s6_sel: begin
                              m4_nxt_st[48:0] = m4_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m4_latch_cmd = m4_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m4_s6_cmd_cur = m4_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m4_s6_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S6_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s7_sel: begin
                              m4_nxt_st[48:0] = m4_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m4_latch_cmd = m4_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m4_s7_cmd_cur = m4_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m4_s7_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S7_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s8_sel: begin
                              m4_nxt_st[48:0] = m4_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m4_latch_cmd = m4_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m4_s8_cmd_cur = m4_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m4_s8_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S8_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s9_sel: begin
                              m4_nxt_st[48:0] = m4_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m4_latch_cmd = m4_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m4_s9_cmd_cur = m4_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m4_s9_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S9_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s10_sel: begin
                              m4_nxt_st[48:0] = m4_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m4_latch_cmd = m4_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m4_s10_cmd_cur = m4_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m4_s10_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S10_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s11_sel: begin
                              m4_nxt_st[48:0] = m4_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m4_latch_cmd = m4_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m4_s11_cmd_cur = m4_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m4_s11_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S11_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             default: begin
                             m4_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m4_nxt_st[48:0] = S_S4_DATA;
end
  S_S5_CMD: begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = s5_hready ? 1'b1 : 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       m4_nxt_st[48:0] = s5_hready  ? S_S5_DATA : S_S5_CMD;
  end
  S_S5_DATA:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b1;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       if(s5_hready)
         begin
           case(1'b1)
             m4_s0_sel: begin
                              m4_nxt_st[48:0] = m4_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m4_latch_cmd = m4_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m4_s0_cmd_cur = m4_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m4_s0_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S0_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s1_sel: begin
                              m4_nxt_st[48:0] = m4_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m4_latch_cmd = m4_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m4_s1_cmd_cur = m4_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m4_s1_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S1_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s2_sel: begin
                              m4_nxt_st[48:0] = m4_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m4_latch_cmd = m4_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m4_s2_cmd_cur = m4_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m4_s2_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S2_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s3_sel: begin
                              m4_nxt_st[48:0] = m4_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m4_latch_cmd = m4_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m4_s3_cmd_cur = m4_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m4_s3_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S3_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s4_sel: begin
                              m4_nxt_st[48:0] = m4_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m4_latch_cmd = m4_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m4_s4_cmd_cur = m4_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m4_s4_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S4_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s5_sel: begin
                              m4_nxt_st[48:0] = S_S5_DATA;
                              m4_s5_cmd_cur = 1'b1;
                             end
             m4_s5_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S5_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s6_sel: begin
                              m4_nxt_st[48:0] = m4_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m4_latch_cmd = m4_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m4_s6_cmd_cur = m4_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m4_s6_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S6_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s7_sel: begin
                              m4_nxt_st[48:0] = m4_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m4_latch_cmd = m4_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m4_s7_cmd_cur = m4_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m4_s7_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S7_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s8_sel: begin
                              m4_nxt_st[48:0] = m4_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m4_latch_cmd = m4_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m4_s8_cmd_cur = m4_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m4_s8_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S8_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s9_sel: begin
                              m4_nxt_st[48:0] = m4_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m4_latch_cmd = m4_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m4_s9_cmd_cur = m4_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m4_s9_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S9_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s10_sel: begin
                              m4_nxt_st[48:0] = m4_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m4_latch_cmd = m4_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m4_s10_cmd_cur = m4_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m4_s10_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S10_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s11_sel: begin
                              m4_nxt_st[48:0] = m4_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m4_latch_cmd = m4_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m4_s11_cmd_cur = m4_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m4_s11_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S11_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             default: begin
                             m4_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m4_nxt_st[48:0] = S_S5_DATA;
end
  S_S6_CMD: begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = s6_hready ? 1'b1 : 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       m4_nxt_st[48:0] = s6_hready  ? S_S6_DATA : S_S6_CMD;
  end
  S_S6_DATA:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b1;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       if(s6_hready)
         begin
           case(1'b1)
             m4_s0_sel: begin
                              m4_nxt_st[48:0] = m4_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m4_latch_cmd = m4_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m4_s0_cmd_cur = m4_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m4_s0_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S0_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s1_sel: begin
                              m4_nxt_st[48:0] = m4_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m4_latch_cmd = m4_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m4_s1_cmd_cur = m4_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m4_s1_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S1_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s2_sel: begin
                              m4_nxt_st[48:0] = m4_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m4_latch_cmd = m4_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m4_s2_cmd_cur = m4_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m4_s2_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S2_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s3_sel: begin
                              m4_nxt_st[48:0] = m4_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m4_latch_cmd = m4_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m4_s3_cmd_cur = m4_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m4_s3_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S3_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s4_sel: begin
                              m4_nxt_st[48:0] = m4_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m4_latch_cmd = m4_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m4_s4_cmd_cur = m4_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m4_s4_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S4_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s5_sel: begin
                              m4_nxt_st[48:0] = m4_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m4_latch_cmd = m4_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m4_s5_cmd_cur = m4_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m4_s5_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S5_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s6_sel: begin
                              m4_nxt_st[48:0] = S_S6_DATA;
                              m4_s6_cmd_cur = 1'b1;
                             end
             m4_s6_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S6_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s7_sel: begin
                              m4_nxt_st[48:0] = m4_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m4_latch_cmd = m4_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m4_s7_cmd_cur = m4_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m4_s7_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S7_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s8_sel: begin
                              m4_nxt_st[48:0] = m4_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m4_latch_cmd = m4_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m4_s8_cmd_cur = m4_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m4_s8_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S8_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s9_sel: begin
                              m4_nxt_st[48:0] = m4_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m4_latch_cmd = m4_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m4_s9_cmd_cur = m4_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m4_s9_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S9_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s10_sel: begin
                              m4_nxt_st[48:0] = m4_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m4_latch_cmd = m4_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m4_s10_cmd_cur = m4_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m4_s10_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S10_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s11_sel: begin
                              m4_nxt_st[48:0] = m4_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m4_latch_cmd = m4_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m4_s11_cmd_cur = m4_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m4_s11_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S11_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             default: begin
                             m4_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m4_nxt_st[48:0] = S_S6_DATA;
end
  S_S7_CMD: begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = s7_hready ? 1'b1 : 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       m4_nxt_st[48:0] = s7_hready  ? S_S7_DATA : S_S7_CMD;
  end
  S_S7_DATA:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b1;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       if(s7_hready)
         begin
           case(1'b1)
             m4_s0_sel: begin
                              m4_nxt_st[48:0] = m4_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m4_latch_cmd = m4_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m4_s0_cmd_cur = m4_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m4_s0_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S0_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s1_sel: begin
                              m4_nxt_st[48:0] = m4_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m4_latch_cmd = m4_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m4_s1_cmd_cur = m4_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m4_s1_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S1_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s2_sel: begin
                              m4_nxt_st[48:0] = m4_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m4_latch_cmd = m4_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m4_s2_cmd_cur = m4_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m4_s2_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S2_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s3_sel: begin
                              m4_nxt_st[48:0] = m4_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m4_latch_cmd = m4_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m4_s3_cmd_cur = m4_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m4_s3_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S3_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s4_sel: begin
                              m4_nxt_st[48:0] = m4_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m4_latch_cmd = m4_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m4_s4_cmd_cur = m4_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m4_s4_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S4_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s5_sel: begin
                              m4_nxt_st[48:0] = m4_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m4_latch_cmd = m4_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m4_s5_cmd_cur = m4_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m4_s5_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S5_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s6_sel: begin
                              m4_nxt_st[48:0] = m4_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m4_latch_cmd = m4_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m4_s6_cmd_cur = m4_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m4_s6_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S6_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s7_sel: begin
                              m4_nxt_st[48:0] = S_S7_DATA;
                              m4_s7_cmd_cur = 1'b1;
                             end
             m4_s7_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S7_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s8_sel: begin
                              m4_nxt_st[48:0] = m4_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m4_latch_cmd = m4_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m4_s8_cmd_cur = m4_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m4_s8_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S8_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s9_sel: begin
                              m4_nxt_st[48:0] = m4_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m4_latch_cmd = m4_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m4_s9_cmd_cur = m4_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m4_s9_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S9_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s10_sel: begin
                              m4_nxt_st[48:0] = m4_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m4_latch_cmd = m4_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m4_s10_cmd_cur = m4_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m4_s10_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S10_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s11_sel: begin
                              m4_nxt_st[48:0] = m4_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m4_latch_cmd = m4_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m4_s11_cmd_cur = m4_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m4_s11_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S11_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             default: begin
                             m4_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m4_nxt_st[48:0] = S_S7_DATA;
end
  S_S8_CMD: begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = s8_hready ? 1'b1 : 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       m4_nxt_st[48:0] = s8_hready  ? S_S8_DATA : S_S8_CMD;
  end
  S_S8_DATA:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b1;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       if(s8_hready)
         begin
           case(1'b1)
             m4_s0_sel: begin
                              m4_nxt_st[48:0] = m4_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m4_latch_cmd = m4_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m4_s0_cmd_cur = m4_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m4_s0_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S0_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s1_sel: begin
                              m4_nxt_st[48:0] = m4_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m4_latch_cmd = m4_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m4_s1_cmd_cur = m4_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m4_s1_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S1_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s2_sel: begin
                              m4_nxt_st[48:0] = m4_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m4_latch_cmd = m4_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m4_s2_cmd_cur = m4_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m4_s2_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S2_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s3_sel: begin
                              m4_nxt_st[48:0] = m4_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m4_latch_cmd = m4_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m4_s3_cmd_cur = m4_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m4_s3_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S3_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s4_sel: begin
                              m4_nxt_st[48:0] = m4_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m4_latch_cmd = m4_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m4_s4_cmd_cur = m4_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m4_s4_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S4_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s5_sel: begin
                              m4_nxt_st[48:0] = m4_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m4_latch_cmd = m4_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m4_s5_cmd_cur = m4_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m4_s5_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S5_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s6_sel: begin
                              m4_nxt_st[48:0] = m4_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m4_latch_cmd = m4_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m4_s6_cmd_cur = m4_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m4_s6_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S6_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s7_sel: begin
                              m4_nxt_st[48:0] = m4_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m4_latch_cmd = m4_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m4_s7_cmd_cur = m4_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m4_s7_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S7_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s8_sel: begin
                              m4_nxt_st[48:0] = S_S8_DATA;
                              m4_s8_cmd_cur = 1'b1;
                             end
             m4_s8_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S8_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s9_sel: begin
                              m4_nxt_st[48:0] = m4_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m4_latch_cmd = m4_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m4_s9_cmd_cur = m4_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m4_s9_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S9_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s10_sel: begin
                              m4_nxt_st[48:0] = m4_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m4_latch_cmd = m4_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m4_s10_cmd_cur = m4_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m4_s10_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S10_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s11_sel: begin
                              m4_nxt_st[48:0] = m4_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m4_latch_cmd = m4_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m4_s11_cmd_cur = m4_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m4_s11_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S11_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             default: begin
                             m4_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m4_nxt_st[48:0] = S_S8_DATA;
end
  S_S9_CMD: begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = s9_hready ? 1'b1 : 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       m4_nxt_st[48:0] = s9_hready  ? S_S9_DATA : S_S9_CMD;
  end
  S_S9_DATA:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b1;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       if(s9_hready)
         begin
           case(1'b1)
             m4_s0_sel: begin
                              m4_nxt_st[48:0] = m4_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m4_latch_cmd = m4_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m4_s0_cmd_cur = m4_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m4_s0_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S0_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s1_sel: begin
                              m4_nxt_st[48:0] = m4_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m4_latch_cmd = m4_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m4_s1_cmd_cur = m4_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m4_s1_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S1_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s2_sel: begin
                              m4_nxt_st[48:0] = m4_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m4_latch_cmd = m4_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m4_s2_cmd_cur = m4_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m4_s2_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S2_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s3_sel: begin
                              m4_nxt_st[48:0] = m4_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m4_latch_cmd = m4_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m4_s3_cmd_cur = m4_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m4_s3_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S3_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s4_sel: begin
                              m4_nxt_st[48:0] = m4_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m4_latch_cmd = m4_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m4_s4_cmd_cur = m4_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m4_s4_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S4_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s5_sel: begin
                              m4_nxt_st[48:0] = m4_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m4_latch_cmd = m4_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m4_s5_cmd_cur = m4_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m4_s5_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S5_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s6_sel: begin
                              m4_nxt_st[48:0] = m4_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m4_latch_cmd = m4_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m4_s6_cmd_cur = m4_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m4_s6_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S6_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s7_sel: begin
                              m4_nxt_st[48:0] = m4_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m4_latch_cmd = m4_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m4_s7_cmd_cur = m4_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m4_s7_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S7_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s8_sel: begin
                              m4_nxt_st[48:0] = m4_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m4_latch_cmd = m4_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m4_s8_cmd_cur = m4_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m4_s8_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S8_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s9_sel: begin
                              m4_nxt_st[48:0] = S_S9_DATA;
                              m4_s9_cmd_cur = 1'b1;
                             end
             m4_s9_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S9_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s10_sel: begin
                              m4_nxt_st[48:0] = m4_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m4_latch_cmd = m4_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m4_s10_cmd_cur = m4_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m4_s10_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S10_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s11_sel: begin
                              m4_nxt_st[48:0] = m4_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m4_latch_cmd = m4_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m4_s11_cmd_cur = m4_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m4_s11_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S11_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             default: begin
                             m4_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m4_nxt_st[48:0] = S_S9_DATA;
end
  S_S10_CMD: begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = s10_hready ? 1'b1 : 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       m4_nxt_st[48:0] = s10_hready  ? S_S10_DATA : S_S10_CMD;
  end
  S_S10_DATA:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b1;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       if(s10_hready)
         begin
           case(1'b1)
             m4_s0_sel: begin
                              m4_nxt_st[48:0] = m4_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m4_latch_cmd = m4_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m4_s0_cmd_cur = m4_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m4_s0_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S0_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s1_sel: begin
                              m4_nxt_st[48:0] = m4_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m4_latch_cmd = m4_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m4_s1_cmd_cur = m4_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m4_s1_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S1_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s2_sel: begin
                              m4_nxt_st[48:0] = m4_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m4_latch_cmd = m4_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m4_s2_cmd_cur = m4_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m4_s2_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S2_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s3_sel: begin
                              m4_nxt_st[48:0] = m4_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m4_latch_cmd = m4_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m4_s3_cmd_cur = m4_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m4_s3_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S3_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s4_sel: begin
                              m4_nxt_st[48:0] = m4_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m4_latch_cmd = m4_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m4_s4_cmd_cur = m4_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m4_s4_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S4_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s5_sel: begin
                              m4_nxt_st[48:0] = m4_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m4_latch_cmd = m4_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m4_s5_cmd_cur = m4_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m4_s5_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S5_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s6_sel: begin
                              m4_nxt_st[48:0] = m4_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m4_latch_cmd = m4_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m4_s6_cmd_cur = m4_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m4_s6_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S6_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s7_sel: begin
                              m4_nxt_st[48:0] = m4_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m4_latch_cmd = m4_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m4_s7_cmd_cur = m4_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m4_s7_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S7_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s8_sel: begin
                              m4_nxt_st[48:0] = m4_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m4_latch_cmd = m4_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m4_s8_cmd_cur = m4_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m4_s8_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S8_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s9_sel: begin
                              m4_nxt_st[48:0] = m4_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m4_latch_cmd = m4_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m4_s9_cmd_cur = m4_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m4_s9_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S9_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s10_sel: begin
                              m4_nxt_st[48:0] = S_S10_DATA;
                              m4_s10_cmd_cur = 1'b1;
                             end
             m4_s10_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S10_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s11_sel: begin
                              m4_nxt_st[48:0] = m4_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m4_latch_cmd = m4_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m4_s11_cmd_cur = m4_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m4_s11_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S11_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             default: begin
                             m4_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m4_nxt_st[48:0] = S_S10_DATA;
end
  S_S11_CMD: begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = s11_hready ? 1'b1 : 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b0;
       m4_nxt_st[48:0] = s11_hready  ? S_S11_DATA : S_S11_CMD;
  end
  S_S11_DATA:begin
       m4_latch_cmd = 1'b0;
       m4_s0_cmd_last = 1'b0;
       m4_s0_cmd_cur = 1'b0;
       m4_s0_data = 1'b0;
       m4_s1_cmd_last = 1'b0;
       m4_s1_cmd_cur = 1'b0;
       m4_s1_data = 1'b0;
       m4_s2_cmd_last = 1'b0;
       m4_s2_cmd_cur = 1'b0;
       m4_s2_data = 1'b0;
       m4_s3_cmd_last = 1'b0;
       m4_s3_cmd_cur = 1'b0;
       m4_s3_data = 1'b0;
       m4_s4_cmd_last = 1'b0;
       m4_s4_cmd_cur = 1'b0;
       m4_s4_data = 1'b0;
       m4_s5_cmd_last = 1'b0;
       m4_s5_cmd_cur = 1'b0;
       m4_s5_data = 1'b0;
       m4_s6_cmd_last = 1'b0;
       m4_s6_cmd_cur = 1'b0;
       m4_s6_data = 1'b0;
       m4_s7_cmd_last = 1'b0;
       m4_s7_cmd_cur = 1'b0;
       m4_s7_data = 1'b0;
       m4_s8_cmd_last = 1'b0;
       m4_s8_cmd_cur = 1'b0;
       m4_s8_data = 1'b0;
       m4_s9_cmd_last = 1'b0;
       m4_s9_cmd_cur = 1'b0;
       m4_s9_data = 1'b0;
       m4_s10_cmd_last = 1'b0;
       m4_s10_cmd_cur = 1'b0;
       m4_s10_data = 1'b0;
       m4_s11_cmd_last = 1'b0;
       m4_s11_cmd_cur = 1'b0;
       m4_s11_data = 1'b1;
       if(s11_hready)
         begin
           case(1'b1)
             m4_s0_sel: begin
                              m4_nxt_st[48:0] = m4_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m4_latch_cmd = m4_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m4_s0_cmd_cur = m4_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m4_s0_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S0_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s1_sel: begin
                              m4_nxt_st[48:0] = m4_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m4_latch_cmd = m4_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m4_s1_cmd_cur = m4_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m4_s1_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S1_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s2_sel: begin
                              m4_nxt_st[48:0] = m4_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m4_latch_cmd = m4_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m4_s2_cmd_cur = m4_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m4_s2_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S2_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s3_sel: begin
                              m4_nxt_st[48:0] = m4_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m4_latch_cmd = m4_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m4_s3_cmd_cur = m4_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m4_s3_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S3_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s4_sel: begin
                              m4_nxt_st[48:0] = m4_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m4_latch_cmd = m4_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m4_s4_cmd_cur = m4_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m4_s4_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S4_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s5_sel: begin
                              m4_nxt_st[48:0] = m4_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m4_latch_cmd = m4_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m4_s5_cmd_cur = m4_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m4_s5_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S5_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s6_sel: begin
                              m4_nxt_st[48:0] = m4_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m4_latch_cmd = m4_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m4_s6_cmd_cur = m4_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m4_s6_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S6_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s7_sel: begin
                              m4_nxt_st[48:0] = m4_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m4_latch_cmd = m4_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m4_s7_cmd_cur = m4_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m4_s7_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S7_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s8_sel: begin
                              m4_nxt_st[48:0] = m4_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m4_latch_cmd = m4_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m4_s8_cmd_cur = m4_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m4_s8_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S8_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s9_sel: begin
                              m4_nxt_st[48:0] = m4_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m4_latch_cmd = m4_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m4_s9_cmd_cur = m4_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m4_s9_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S9_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s10_sel: begin
                              m4_nxt_st[48:0] = m4_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m4_latch_cmd = m4_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m4_s10_cmd_cur = m4_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m4_s10_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S10_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             m4_s11_sel: begin
                              m4_nxt_st[48:0] = S_S11_DATA;
                              m4_s11_cmd_cur = 1'b1;
                             end
             m4_s11_wt_sel: begin
                                 m4_nxt_st[48:0] = S_S11_GNT;
                                 m4_latch_cmd = 1'b1;
                               end
             default: begin
                             m4_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m4_nxt_st[48:0] = S_S11_DATA;
end
  default: begin
             m4_latch_cmd = 1'b0;
             m4_s0_cmd_last = 1'b0;
             m4_s0_cmd_cur = 1'b0;
             m4_s0_data = 1'b0;
             m4_s1_cmd_last = 1'b0;
             m4_s1_cmd_cur = 1'b0;
             m4_s1_data = 1'b0;
             m4_s2_cmd_last = 1'b0;
             m4_s2_cmd_cur = 1'b0;
             m4_s2_data = 1'b0;
             m4_s3_cmd_last = 1'b0;
             m4_s3_cmd_cur = 1'b0;
             m4_s3_data = 1'b0;
             m4_s4_cmd_last = 1'b0;
             m4_s4_cmd_cur = 1'b0;
             m4_s4_data = 1'b0;
             m4_s5_cmd_last = 1'b0;
             m4_s5_cmd_cur = 1'b0;
             m4_s5_data = 1'b0;
             m4_s6_cmd_last = 1'b0;
             m4_s6_cmd_cur = 1'b0;
             m4_s6_data = 1'b0;
             m4_s7_cmd_last = 1'b0;
             m4_s7_cmd_cur = 1'b0;
             m4_s7_data = 1'b0;
             m4_s8_cmd_last = 1'b0;
             m4_s8_cmd_cur = 1'b0;
             m4_s8_data = 1'b0;
             m4_s9_cmd_last = 1'b0;
             m4_s9_cmd_cur = 1'b0;
             m4_s9_data = 1'b0;
             m4_s10_cmd_last = 1'b0;
             m4_s10_cmd_cur = 1'b0;
             m4_s10_data = 1'b0;
             m4_s11_cmd_last = 1'b0;
             m4_s11_cmd_cur = 1'b0;
             m4_s11_data = 1'b0;
             m4_nxt_st[48:0] = S_IDLE;
  end
endcase
end
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
       m5_cur_st[48:0] <= S_IDLE;
    else
       m5_cur_st[48:0] <= m5_nxt_st[48:0];
  end
always @ (*)
begin
case(m5_cur_st[48:0])
  S_IDLE:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       case(1'b1)
         m5_s0_sel: begin
                          m5_nxt_st[48:0] = m5_s0_hld ? S_S0_WAIT : (s0_hready ? S_S0_DATA : S_S0_CMD);
                          m5_latch_cmd = m5_s0_hld ? 1'b1 : (s0_hready ? 1'b0 : 1'b1);
                          m5_s0_cmd_cur = m5_s0_hld ? 1'b0 : (s0_hready ? 1'b1 : 1'b0);
                        end
         m5_s0_wt_sel: begin
                             m5_nxt_st[48:0] = S_S0_GNT;
                             m5_latch_cmd = 1'b1;
                           end
         m5_s1_sel: begin
                          m5_nxt_st[48:0] = m5_s1_hld ? S_S1_WAIT : (s1_hready ? S_S1_DATA : S_S1_CMD);
                          m5_latch_cmd = m5_s1_hld ? 1'b1 : (s1_hready ? 1'b0 : 1'b1);
                          m5_s1_cmd_cur = m5_s1_hld ? 1'b0 : (s1_hready ? 1'b1 : 1'b0);
                        end
         m5_s1_wt_sel: begin
                             m5_nxt_st[48:0] = S_S1_GNT;
                             m5_latch_cmd = 1'b1;
                           end
         m5_s2_sel: begin
                          m5_nxt_st[48:0] = m5_s2_hld ? S_S2_WAIT : (s2_hready ? S_S2_DATA : S_S2_CMD);
                          m5_latch_cmd = m5_s2_hld ? 1'b1 : (s2_hready ? 1'b0 : 1'b1);
                          m5_s2_cmd_cur = m5_s2_hld ? 1'b0 : (s2_hready ? 1'b1 : 1'b0);
                        end
         m5_s2_wt_sel: begin
                             m5_nxt_st[48:0] = S_S2_GNT;
                             m5_latch_cmd = 1'b1;
                           end
         m5_s3_sel: begin
                          m5_nxt_st[48:0] = m5_s3_hld ? S_S3_WAIT : (s3_hready ? S_S3_DATA : S_S3_CMD);
                          m5_latch_cmd = m5_s3_hld ? 1'b1 : (s3_hready ? 1'b0 : 1'b1);
                          m5_s3_cmd_cur = m5_s3_hld ? 1'b0 : (s3_hready ? 1'b1 : 1'b0);
                        end
         m5_s3_wt_sel: begin
                             m5_nxt_st[48:0] = S_S3_GNT;
                             m5_latch_cmd = 1'b1;
                           end
         m5_s4_sel: begin
                          m5_nxt_st[48:0] = m5_s4_hld ? S_S4_WAIT : (s4_hready ? S_S4_DATA : S_S4_CMD);
                          m5_latch_cmd = m5_s4_hld ? 1'b1 : (s4_hready ? 1'b0 : 1'b1);
                          m5_s4_cmd_cur = m5_s4_hld ? 1'b0 : (s4_hready ? 1'b1 : 1'b0);
                        end
         m5_s4_wt_sel: begin
                             m5_nxt_st[48:0] = S_S4_GNT;
                             m5_latch_cmd = 1'b1;
                           end
         m5_s5_sel: begin
                          m5_nxt_st[48:0] = m5_s5_hld ? S_S5_WAIT : (s5_hready ? S_S5_DATA : S_S5_CMD);
                          m5_latch_cmd = m5_s5_hld ? 1'b1 : (s5_hready ? 1'b0 : 1'b1);
                          m5_s5_cmd_cur = m5_s5_hld ? 1'b0 : (s5_hready ? 1'b1 : 1'b0);
                        end
         m5_s5_wt_sel: begin
                             m5_nxt_st[48:0] = S_S5_GNT;
                             m5_latch_cmd = 1'b1;
                           end
         m5_s6_sel: begin
                          m5_nxt_st[48:0] = m5_s6_hld ? S_S6_WAIT : (s6_hready ? S_S6_DATA : S_S6_CMD);
                          m5_latch_cmd = m5_s6_hld ? 1'b1 : (s6_hready ? 1'b0 : 1'b1);
                          m5_s6_cmd_cur = m5_s6_hld ? 1'b0 : (s6_hready ? 1'b1 : 1'b0);
                        end
         m5_s6_wt_sel: begin
                             m5_nxt_st[48:0] = S_S6_GNT;
                             m5_latch_cmd = 1'b1;
                           end
         m5_s7_sel: begin
                          m5_nxt_st[48:0] = m5_s7_hld ? S_S7_WAIT : (s7_hready ? S_S7_DATA : S_S7_CMD);
                          m5_latch_cmd = m5_s7_hld ? 1'b1 : (s7_hready ? 1'b0 : 1'b1);
                          m5_s7_cmd_cur = m5_s7_hld ? 1'b0 : (s7_hready ? 1'b1 : 1'b0);
                        end
         m5_s7_wt_sel: begin
                             m5_nxt_st[48:0] = S_S7_GNT;
                             m5_latch_cmd = 1'b1;
                           end
         m5_s8_sel: begin
                          m5_nxt_st[48:0] = m5_s8_hld ? S_S8_WAIT : (s8_hready ? S_S8_DATA : S_S8_CMD);
                          m5_latch_cmd = m5_s8_hld ? 1'b1 : (s8_hready ? 1'b0 : 1'b1);
                          m5_s8_cmd_cur = m5_s8_hld ? 1'b0 : (s8_hready ? 1'b1 : 1'b0);
                        end
         m5_s8_wt_sel: begin
                             m5_nxt_st[48:0] = S_S8_GNT;
                             m5_latch_cmd = 1'b1;
                           end
         m5_s9_sel: begin
                          m5_nxt_st[48:0] = m5_s9_hld ? S_S9_WAIT : (s9_hready ? S_S9_DATA : S_S9_CMD);
                          m5_latch_cmd = m5_s9_hld ? 1'b1 : (s9_hready ? 1'b0 : 1'b1);
                          m5_s9_cmd_cur = m5_s9_hld ? 1'b0 : (s9_hready ? 1'b1 : 1'b0);
                        end
         m5_s9_wt_sel: begin
                             m5_nxt_st[48:0] = S_S9_GNT;
                             m5_latch_cmd = 1'b1;
                           end
         m5_s10_sel: begin
                          m5_nxt_st[48:0] = m5_s10_hld ? S_S10_WAIT : (s10_hready ? S_S10_DATA : S_S10_CMD);
                          m5_latch_cmd = m5_s10_hld ? 1'b1 : (s10_hready ? 1'b0 : 1'b1);
                          m5_s10_cmd_cur = m5_s10_hld ? 1'b0 : (s10_hready ? 1'b1 : 1'b0);
                        end
         m5_s10_wt_sel: begin
                             m5_nxt_st[48:0] = S_S10_GNT;
                             m5_latch_cmd = 1'b1;
                           end
         m5_s11_sel: begin
                          m5_nxt_st[48:0] = m5_s11_hld ? S_S11_WAIT : (s11_hready ? S_S11_DATA : S_S11_CMD);
                          m5_latch_cmd = m5_s11_hld ? 1'b1 : (s11_hready ? 1'b0 : 1'b1);
                          m5_s11_cmd_cur = m5_s11_hld ? 1'b0 : (s11_hready ? 1'b1 : 1'b0);
                        end
         m5_s11_wt_sel: begin
                             m5_nxt_st[48:0] = S_S11_GNT;
                             m5_latch_cmd = 1'b1;
                           end
         default: begin
                          m5_nxt_st[48:0] = S_IDLE;
                  end
       endcase
  end
  S_S0_GNT:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       case(1'b1)
         m5_s0_sel: begin
                          m5_nxt_st[48:0] = m5_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                          m5_s0_cmd_last = m5_s0_hld ? 1'b0 : (s0_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m5_nxt_st[48:0] = S_S0_GNT;
                  end
       endcase
  end
  S_S1_GNT:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       case(1'b1)
         m5_s1_sel: begin
                          m5_nxt_st[48:0] = m5_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                          m5_s1_cmd_last = m5_s1_hld ? 1'b0 : (s1_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m5_nxt_st[48:0] = S_S1_GNT;
                  end
       endcase
  end
  S_S2_GNT:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       case(1'b1)
         m5_s2_sel: begin
                          m5_nxt_st[48:0] = m5_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                          m5_s2_cmd_last = m5_s2_hld ? 1'b0 : (s2_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m5_nxt_st[48:0] = S_S2_GNT;
                  end
       endcase
  end
  S_S3_GNT:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       case(1'b1)
         m5_s3_sel: begin
                          m5_nxt_st[48:0] = m5_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                          m5_s3_cmd_last = m5_s3_hld ? 1'b0 : (s3_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m5_nxt_st[48:0] = S_S3_GNT;
                  end
       endcase
  end
  S_S4_GNT:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       case(1'b1)
         m5_s4_sel: begin
                          m5_nxt_st[48:0] = m5_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                          m5_s4_cmd_last = m5_s4_hld ? 1'b0 : (s4_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m5_nxt_st[48:0] = S_S4_GNT;
                  end
       endcase
  end
  S_S5_GNT:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       case(1'b1)
         m5_s5_sel: begin
                          m5_nxt_st[48:0] = m5_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                          m5_s5_cmd_last = m5_s5_hld ? 1'b0 : (s5_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m5_nxt_st[48:0] = S_S5_GNT;
                  end
       endcase
  end
  S_S6_GNT:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       case(1'b1)
         m5_s6_sel: begin
                          m5_nxt_st[48:0] = m5_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                          m5_s6_cmd_last = m5_s6_hld ? 1'b0 : (s6_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m5_nxt_st[48:0] = S_S6_GNT;
                  end
       endcase
  end
  S_S7_GNT:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       case(1'b1)
         m5_s7_sel: begin
                          m5_nxt_st[48:0] = m5_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                          m5_s7_cmd_last = m5_s7_hld ? 1'b0 : (s7_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m5_nxt_st[48:0] = S_S7_GNT;
                  end
       endcase
  end
  S_S8_GNT:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       case(1'b1)
         m5_s8_sel: begin
                          m5_nxt_st[48:0] = m5_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                          m5_s8_cmd_last = m5_s8_hld ? 1'b0 : (s8_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m5_nxt_st[48:0] = S_S8_GNT;
                  end
       endcase
  end
  S_S9_GNT:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       case(1'b1)
         m5_s9_sel: begin
                          m5_nxt_st[48:0] = m5_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                          m5_s9_cmd_last = m5_s9_hld ? 1'b0 : (s9_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m5_nxt_st[48:0] = S_S9_GNT;
                  end
       endcase
  end
  S_S10_GNT:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       case(1'b1)
         m5_s10_sel: begin
                          m5_nxt_st[48:0] = m5_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                          m5_s10_cmd_last = m5_s10_hld ? 1'b0 : (s10_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m5_nxt_st[48:0] = S_S10_GNT;
                  end
       endcase
  end
  S_S11_GNT:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       case(1'b1)
         m5_s11_sel: begin
                          m5_nxt_st[48:0] = m5_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                          m5_s11_cmd_last = m5_s11_hld ? 1'b0 : (s11_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m5_nxt_st[48:0] = S_S11_GNT;
                  end
       endcase
  end
  S_S0_WAIT:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       case(1'b1)
         ~m5_s0_hld: begin
                          m5_nxt_st[48:0] = m5_s0_wt_sel ? S_S0_GNT : s0_hready ? S_S0_DATA : S_S0_CMD;
                          m5_s0_cmd_last = m5_s0_wt_sel ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m5_nxt_st[48:0] = S_S0_WAIT;
                  end
       endcase
  end
  S_S1_WAIT:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       case(1'b1)
         ~m5_s1_hld: begin
                          m5_nxt_st[48:0] = m5_s1_wt_sel ? S_S1_GNT : s1_hready ? S_S1_DATA : S_S1_CMD;
                          m5_s1_cmd_last = m5_s1_wt_sel ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m5_nxt_st[48:0] = S_S1_WAIT;
                  end
       endcase
  end
  S_S2_WAIT:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       case(1'b1)
         ~m5_s2_hld: begin
                          m5_nxt_st[48:0] = m5_s2_wt_sel ? S_S2_GNT : s2_hready ? S_S2_DATA : S_S2_CMD;
                          m5_s2_cmd_last = m5_s2_wt_sel ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m5_nxt_st[48:0] = S_S2_WAIT;
                  end
       endcase
  end
  S_S3_WAIT:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       case(1'b1)
         ~m5_s3_hld: begin
                          m5_nxt_st[48:0] = m5_s3_wt_sel ? S_S3_GNT : s3_hready ? S_S3_DATA : S_S3_CMD;
                          m5_s3_cmd_last = m5_s3_wt_sel ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m5_nxt_st[48:0] = S_S3_WAIT;
                  end
       endcase
  end
  S_S4_WAIT:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       case(1'b1)
         ~m5_s4_hld: begin
                          m5_nxt_st[48:0] = m5_s4_wt_sel ? S_S4_GNT : s4_hready ? S_S4_DATA : S_S4_CMD;
                          m5_s4_cmd_last = m5_s4_wt_sel ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m5_nxt_st[48:0] = S_S4_WAIT;
                  end
       endcase
  end
  S_S5_WAIT:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       case(1'b1)
         ~m5_s5_hld: begin
                          m5_nxt_st[48:0] = m5_s5_wt_sel ? S_S5_GNT : s5_hready ? S_S5_DATA : S_S5_CMD;
                          m5_s5_cmd_last = m5_s5_wt_sel ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m5_nxt_st[48:0] = S_S5_WAIT;
                  end
       endcase
  end
  S_S6_WAIT:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       case(1'b1)
         ~m5_s6_hld: begin
                          m5_nxt_st[48:0] = m5_s6_wt_sel ? S_S6_GNT : s6_hready ? S_S6_DATA : S_S6_CMD;
                          m5_s6_cmd_last = m5_s6_wt_sel ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m5_nxt_st[48:0] = S_S6_WAIT;
                  end
       endcase
  end
  S_S7_WAIT:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       case(1'b1)
         ~m5_s7_hld: begin
                          m5_nxt_st[48:0] = m5_s7_wt_sel ? S_S7_GNT : s7_hready ? S_S7_DATA : S_S7_CMD;
                          m5_s7_cmd_last = m5_s7_wt_sel ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m5_nxt_st[48:0] = S_S7_WAIT;
                  end
       endcase
  end
  S_S8_WAIT:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       case(1'b1)
         ~m5_s8_hld: begin
                          m5_nxt_st[48:0] = m5_s8_wt_sel ? S_S8_GNT : s8_hready ? S_S8_DATA : S_S8_CMD;
                          m5_s8_cmd_last = m5_s8_wt_sel ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m5_nxt_st[48:0] = S_S8_WAIT;
                  end
       endcase
  end
  S_S9_WAIT:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       case(1'b1)
         ~m5_s9_hld: begin
                          m5_nxt_st[48:0] = m5_s9_wt_sel ? S_S9_GNT : s9_hready ? S_S9_DATA : S_S9_CMD;
                          m5_s9_cmd_last = m5_s9_wt_sel ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m5_nxt_st[48:0] = S_S9_WAIT;
                  end
       endcase
  end
  S_S10_WAIT:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       case(1'b1)
         ~m5_s10_hld: begin
                          m5_nxt_st[48:0] = m5_s10_wt_sel ? S_S10_GNT : s10_hready ? S_S10_DATA : S_S10_CMD;
                          m5_s10_cmd_last = m5_s10_wt_sel ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m5_nxt_st[48:0] = S_S10_WAIT;
                  end
       endcase
  end
  S_S11_WAIT:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       case(1'b1)
         ~m5_s11_hld: begin
                          m5_nxt_st[48:0] = m5_s11_wt_sel ? S_S11_GNT : s11_hready ? S_S11_DATA : S_S11_CMD;
                          m5_s11_cmd_last = m5_s11_wt_sel ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m5_nxt_st[48:0] = S_S11_WAIT;
                  end
       endcase
  end
  S_S0_CMD: begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = s0_hready ? 1'b1 : 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       m5_nxt_st[48:0] = s0_hready  ? S_S0_DATA : S_S0_CMD;
  end
  S_S0_DATA:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b1;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       if(s0_hready)
         begin
           case(1'b1)
             m5_s0_sel: begin
                              m5_nxt_st[48:0] = S_S0_DATA;
                              m5_s0_cmd_cur = 1'b1;
                             end
             m5_s0_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S0_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s1_sel: begin
                              m5_nxt_st[48:0] = m5_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m5_latch_cmd = m5_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m5_s1_cmd_cur = m5_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m5_s1_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S1_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s2_sel: begin
                              m5_nxt_st[48:0] = m5_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m5_latch_cmd = m5_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m5_s2_cmd_cur = m5_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m5_s2_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S2_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s3_sel: begin
                              m5_nxt_st[48:0] = m5_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m5_latch_cmd = m5_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m5_s3_cmd_cur = m5_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m5_s3_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S3_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s4_sel: begin
                              m5_nxt_st[48:0] = m5_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m5_latch_cmd = m5_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m5_s4_cmd_cur = m5_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m5_s4_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S4_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s5_sel: begin
                              m5_nxt_st[48:0] = m5_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m5_latch_cmd = m5_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m5_s5_cmd_cur = m5_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m5_s5_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S5_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s6_sel: begin
                              m5_nxt_st[48:0] = m5_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m5_latch_cmd = m5_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m5_s6_cmd_cur = m5_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m5_s6_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S6_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s7_sel: begin
                              m5_nxt_st[48:0] = m5_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m5_latch_cmd = m5_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m5_s7_cmd_cur = m5_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m5_s7_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S7_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s8_sel: begin
                              m5_nxt_st[48:0] = m5_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m5_latch_cmd = m5_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m5_s8_cmd_cur = m5_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m5_s8_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S8_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s9_sel: begin
                              m5_nxt_st[48:0] = m5_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m5_latch_cmd = m5_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m5_s9_cmd_cur = m5_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m5_s9_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S9_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s10_sel: begin
                              m5_nxt_st[48:0] = m5_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m5_latch_cmd = m5_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m5_s10_cmd_cur = m5_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m5_s10_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S10_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s11_sel: begin
                              m5_nxt_st[48:0] = m5_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m5_latch_cmd = m5_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m5_s11_cmd_cur = m5_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m5_s11_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S11_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             default: begin
                             m5_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m5_nxt_st[48:0] = S_S0_DATA;
end
  S_S1_CMD: begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = s1_hready ? 1'b1 : 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       m5_nxt_st[48:0] = s1_hready  ? S_S1_DATA : S_S1_CMD;
  end
  S_S1_DATA:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b1;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       if(s1_hready)
         begin
           case(1'b1)
             m5_s0_sel: begin
                              m5_nxt_st[48:0] = m5_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m5_latch_cmd = m5_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m5_s0_cmd_cur = m5_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m5_s0_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S0_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s1_sel: begin
                              m5_nxt_st[48:0] = S_S1_DATA;
                              m5_s1_cmd_cur = 1'b1;
                             end
             m5_s1_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S1_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s2_sel: begin
                              m5_nxt_st[48:0] = m5_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m5_latch_cmd = m5_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m5_s2_cmd_cur = m5_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m5_s2_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S2_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s3_sel: begin
                              m5_nxt_st[48:0] = m5_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m5_latch_cmd = m5_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m5_s3_cmd_cur = m5_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m5_s3_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S3_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s4_sel: begin
                              m5_nxt_st[48:0] = m5_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m5_latch_cmd = m5_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m5_s4_cmd_cur = m5_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m5_s4_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S4_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s5_sel: begin
                              m5_nxt_st[48:0] = m5_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m5_latch_cmd = m5_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m5_s5_cmd_cur = m5_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m5_s5_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S5_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s6_sel: begin
                              m5_nxt_st[48:0] = m5_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m5_latch_cmd = m5_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m5_s6_cmd_cur = m5_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m5_s6_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S6_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s7_sel: begin
                              m5_nxt_st[48:0] = m5_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m5_latch_cmd = m5_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m5_s7_cmd_cur = m5_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m5_s7_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S7_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s8_sel: begin
                              m5_nxt_st[48:0] = m5_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m5_latch_cmd = m5_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m5_s8_cmd_cur = m5_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m5_s8_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S8_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s9_sel: begin
                              m5_nxt_st[48:0] = m5_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m5_latch_cmd = m5_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m5_s9_cmd_cur = m5_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m5_s9_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S9_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s10_sel: begin
                              m5_nxt_st[48:0] = m5_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m5_latch_cmd = m5_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m5_s10_cmd_cur = m5_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m5_s10_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S10_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s11_sel: begin
                              m5_nxt_st[48:0] = m5_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m5_latch_cmd = m5_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m5_s11_cmd_cur = m5_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m5_s11_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S11_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             default: begin
                             m5_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m5_nxt_st[48:0] = S_S1_DATA;
end
  S_S2_CMD: begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = s2_hready ? 1'b1 : 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       m5_nxt_st[48:0] = s2_hready  ? S_S2_DATA : S_S2_CMD;
  end
  S_S2_DATA:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b1;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       if(s2_hready)
         begin
           case(1'b1)
             m5_s0_sel: begin
                              m5_nxt_st[48:0] = m5_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m5_latch_cmd = m5_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m5_s0_cmd_cur = m5_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m5_s0_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S0_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s1_sel: begin
                              m5_nxt_st[48:0] = m5_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m5_latch_cmd = m5_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m5_s1_cmd_cur = m5_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m5_s1_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S1_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s2_sel: begin
                              m5_nxt_st[48:0] = S_S2_DATA;
                              m5_s2_cmd_cur = 1'b1;
                             end
             m5_s2_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S2_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s3_sel: begin
                              m5_nxt_st[48:0] = m5_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m5_latch_cmd = m5_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m5_s3_cmd_cur = m5_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m5_s3_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S3_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s4_sel: begin
                              m5_nxt_st[48:0] = m5_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m5_latch_cmd = m5_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m5_s4_cmd_cur = m5_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m5_s4_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S4_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s5_sel: begin
                              m5_nxt_st[48:0] = m5_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m5_latch_cmd = m5_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m5_s5_cmd_cur = m5_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m5_s5_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S5_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s6_sel: begin
                              m5_nxt_st[48:0] = m5_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m5_latch_cmd = m5_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m5_s6_cmd_cur = m5_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m5_s6_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S6_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s7_sel: begin
                              m5_nxt_st[48:0] = m5_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m5_latch_cmd = m5_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m5_s7_cmd_cur = m5_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m5_s7_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S7_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s8_sel: begin
                              m5_nxt_st[48:0] = m5_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m5_latch_cmd = m5_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m5_s8_cmd_cur = m5_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m5_s8_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S8_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s9_sel: begin
                              m5_nxt_st[48:0] = m5_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m5_latch_cmd = m5_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m5_s9_cmd_cur = m5_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m5_s9_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S9_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s10_sel: begin
                              m5_nxt_st[48:0] = m5_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m5_latch_cmd = m5_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m5_s10_cmd_cur = m5_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m5_s10_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S10_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s11_sel: begin
                              m5_nxt_st[48:0] = m5_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m5_latch_cmd = m5_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m5_s11_cmd_cur = m5_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m5_s11_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S11_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             default: begin
                             m5_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m5_nxt_st[48:0] = S_S2_DATA;
end
  S_S3_CMD: begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = s3_hready ? 1'b1 : 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       m5_nxt_st[48:0] = s3_hready  ? S_S3_DATA : S_S3_CMD;
  end
  S_S3_DATA:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b1;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       if(s3_hready)
         begin
           case(1'b1)
             m5_s0_sel: begin
                              m5_nxt_st[48:0] = m5_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m5_latch_cmd = m5_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m5_s0_cmd_cur = m5_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m5_s0_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S0_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s1_sel: begin
                              m5_nxt_st[48:0] = m5_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m5_latch_cmd = m5_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m5_s1_cmd_cur = m5_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m5_s1_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S1_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s2_sel: begin
                              m5_nxt_st[48:0] = m5_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m5_latch_cmd = m5_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m5_s2_cmd_cur = m5_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m5_s2_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S2_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s3_sel: begin
                              m5_nxt_st[48:0] = S_S3_DATA;
                              m5_s3_cmd_cur = 1'b1;
                             end
             m5_s3_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S3_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s4_sel: begin
                              m5_nxt_st[48:0] = m5_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m5_latch_cmd = m5_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m5_s4_cmd_cur = m5_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m5_s4_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S4_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s5_sel: begin
                              m5_nxt_st[48:0] = m5_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m5_latch_cmd = m5_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m5_s5_cmd_cur = m5_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m5_s5_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S5_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s6_sel: begin
                              m5_nxt_st[48:0] = m5_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m5_latch_cmd = m5_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m5_s6_cmd_cur = m5_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m5_s6_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S6_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s7_sel: begin
                              m5_nxt_st[48:0] = m5_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m5_latch_cmd = m5_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m5_s7_cmd_cur = m5_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m5_s7_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S7_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s8_sel: begin
                              m5_nxt_st[48:0] = m5_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m5_latch_cmd = m5_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m5_s8_cmd_cur = m5_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m5_s8_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S8_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s9_sel: begin
                              m5_nxt_st[48:0] = m5_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m5_latch_cmd = m5_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m5_s9_cmd_cur = m5_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m5_s9_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S9_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s10_sel: begin
                              m5_nxt_st[48:0] = m5_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m5_latch_cmd = m5_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m5_s10_cmd_cur = m5_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m5_s10_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S10_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s11_sel: begin
                              m5_nxt_st[48:0] = m5_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m5_latch_cmd = m5_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m5_s11_cmd_cur = m5_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m5_s11_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S11_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             default: begin
                             m5_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m5_nxt_st[48:0] = S_S3_DATA;
end
  S_S4_CMD: begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = s4_hready ? 1'b1 : 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       m5_nxt_st[48:0] = s4_hready  ? S_S4_DATA : S_S4_CMD;
  end
  S_S4_DATA:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b1;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       if(s4_hready)
         begin
           case(1'b1)
             m5_s0_sel: begin
                              m5_nxt_st[48:0] = m5_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m5_latch_cmd = m5_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m5_s0_cmd_cur = m5_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m5_s0_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S0_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s1_sel: begin
                              m5_nxt_st[48:0] = m5_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m5_latch_cmd = m5_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m5_s1_cmd_cur = m5_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m5_s1_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S1_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s2_sel: begin
                              m5_nxt_st[48:0] = m5_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m5_latch_cmd = m5_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m5_s2_cmd_cur = m5_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m5_s2_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S2_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s3_sel: begin
                              m5_nxt_st[48:0] = m5_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m5_latch_cmd = m5_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m5_s3_cmd_cur = m5_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m5_s3_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S3_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s4_sel: begin
                              m5_nxt_st[48:0] = S_S4_DATA;
                              m5_s4_cmd_cur = 1'b1;
                             end
             m5_s4_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S4_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s5_sel: begin
                              m5_nxt_st[48:0] = m5_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m5_latch_cmd = m5_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m5_s5_cmd_cur = m5_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m5_s5_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S5_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s6_sel: begin
                              m5_nxt_st[48:0] = m5_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m5_latch_cmd = m5_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m5_s6_cmd_cur = m5_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m5_s6_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S6_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s7_sel: begin
                              m5_nxt_st[48:0] = m5_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m5_latch_cmd = m5_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m5_s7_cmd_cur = m5_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m5_s7_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S7_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s8_sel: begin
                              m5_nxt_st[48:0] = m5_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m5_latch_cmd = m5_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m5_s8_cmd_cur = m5_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m5_s8_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S8_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s9_sel: begin
                              m5_nxt_st[48:0] = m5_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m5_latch_cmd = m5_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m5_s9_cmd_cur = m5_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m5_s9_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S9_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s10_sel: begin
                              m5_nxt_st[48:0] = m5_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m5_latch_cmd = m5_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m5_s10_cmd_cur = m5_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m5_s10_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S10_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s11_sel: begin
                              m5_nxt_st[48:0] = m5_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m5_latch_cmd = m5_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m5_s11_cmd_cur = m5_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m5_s11_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S11_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             default: begin
                             m5_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m5_nxt_st[48:0] = S_S4_DATA;
end
  S_S5_CMD: begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = s5_hready ? 1'b1 : 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       m5_nxt_st[48:0] = s5_hready  ? S_S5_DATA : S_S5_CMD;
  end
  S_S5_DATA:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b1;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       if(s5_hready)
         begin
           case(1'b1)
             m5_s0_sel: begin
                              m5_nxt_st[48:0] = m5_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m5_latch_cmd = m5_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m5_s0_cmd_cur = m5_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m5_s0_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S0_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s1_sel: begin
                              m5_nxt_st[48:0] = m5_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m5_latch_cmd = m5_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m5_s1_cmd_cur = m5_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m5_s1_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S1_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s2_sel: begin
                              m5_nxt_st[48:0] = m5_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m5_latch_cmd = m5_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m5_s2_cmd_cur = m5_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m5_s2_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S2_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s3_sel: begin
                              m5_nxt_st[48:0] = m5_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m5_latch_cmd = m5_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m5_s3_cmd_cur = m5_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m5_s3_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S3_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s4_sel: begin
                              m5_nxt_st[48:0] = m5_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m5_latch_cmd = m5_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m5_s4_cmd_cur = m5_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m5_s4_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S4_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s5_sel: begin
                              m5_nxt_st[48:0] = S_S5_DATA;
                              m5_s5_cmd_cur = 1'b1;
                             end
             m5_s5_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S5_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s6_sel: begin
                              m5_nxt_st[48:0] = m5_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m5_latch_cmd = m5_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m5_s6_cmd_cur = m5_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m5_s6_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S6_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s7_sel: begin
                              m5_nxt_st[48:0] = m5_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m5_latch_cmd = m5_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m5_s7_cmd_cur = m5_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m5_s7_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S7_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s8_sel: begin
                              m5_nxt_st[48:0] = m5_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m5_latch_cmd = m5_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m5_s8_cmd_cur = m5_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m5_s8_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S8_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s9_sel: begin
                              m5_nxt_st[48:0] = m5_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m5_latch_cmd = m5_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m5_s9_cmd_cur = m5_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m5_s9_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S9_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s10_sel: begin
                              m5_nxt_st[48:0] = m5_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m5_latch_cmd = m5_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m5_s10_cmd_cur = m5_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m5_s10_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S10_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s11_sel: begin
                              m5_nxt_st[48:0] = m5_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m5_latch_cmd = m5_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m5_s11_cmd_cur = m5_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m5_s11_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S11_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             default: begin
                             m5_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m5_nxt_st[48:0] = S_S5_DATA;
end
  S_S6_CMD: begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = s6_hready ? 1'b1 : 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       m5_nxt_st[48:0] = s6_hready  ? S_S6_DATA : S_S6_CMD;
  end
  S_S6_DATA:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b1;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       if(s6_hready)
         begin
           case(1'b1)
             m5_s0_sel: begin
                              m5_nxt_st[48:0] = m5_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m5_latch_cmd = m5_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m5_s0_cmd_cur = m5_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m5_s0_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S0_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s1_sel: begin
                              m5_nxt_st[48:0] = m5_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m5_latch_cmd = m5_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m5_s1_cmd_cur = m5_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m5_s1_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S1_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s2_sel: begin
                              m5_nxt_st[48:0] = m5_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m5_latch_cmd = m5_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m5_s2_cmd_cur = m5_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m5_s2_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S2_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s3_sel: begin
                              m5_nxt_st[48:0] = m5_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m5_latch_cmd = m5_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m5_s3_cmd_cur = m5_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m5_s3_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S3_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s4_sel: begin
                              m5_nxt_st[48:0] = m5_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m5_latch_cmd = m5_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m5_s4_cmd_cur = m5_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m5_s4_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S4_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s5_sel: begin
                              m5_nxt_st[48:0] = m5_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m5_latch_cmd = m5_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m5_s5_cmd_cur = m5_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m5_s5_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S5_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s6_sel: begin
                              m5_nxt_st[48:0] = S_S6_DATA;
                              m5_s6_cmd_cur = 1'b1;
                             end
             m5_s6_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S6_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s7_sel: begin
                              m5_nxt_st[48:0] = m5_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m5_latch_cmd = m5_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m5_s7_cmd_cur = m5_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m5_s7_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S7_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s8_sel: begin
                              m5_nxt_st[48:0] = m5_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m5_latch_cmd = m5_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m5_s8_cmd_cur = m5_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m5_s8_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S8_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s9_sel: begin
                              m5_nxt_st[48:0] = m5_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m5_latch_cmd = m5_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m5_s9_cmd_cur = m5_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m5_s9_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S9_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s10_sel: begin
                              m5_nxt_st[48:0] = m5_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m5_latch_cmd = m5_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m5_s10_cmd_cur = m5_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m5_s10_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S10_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s11_sel: begin
                              m5_nxt_st[48:0] = m5_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m5_latch_cmd = m5_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m5_s11_cmd_cur = m5_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m5_s11_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S11_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             default: begin
                             m5_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m5_nxt_st[48:0] = S_S6_DATA;
end
  S_S7_CMD: begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = s7_hready ? 1'b1 : 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       m5_nxt_st[48:0] = s7_hready  ? S_S7_DATA : S_S7_CMD;
  end
  S_S7_DATA:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b1;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       if(s7_hready)
         begin
           case(1'b1)
             m5_s0_sel: begin
                              m5_nxt_st[48:0] = m5_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m5_latch_cmd = m5_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m5_s0_cmd_cur = m5_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m5_s0_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S0_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s1_sel: begin
                              m5_nxt_st[48:0] = m5_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m5_latch_cmd = m5_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m5_s1_cmd_cur = m5_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m5_s1_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S1_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s2_sel: begin
                              m5_nxt_st[48:0] = m5_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m5_latch_cmd = m5_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m5_s2_cmd_cur = m5_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m5_s2_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S2_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s3_sel: begin
                              m5_nxt_st[48:0] = m5_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m5_latch_cmd = m5_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m5_s3_cmd_cur = m5_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m5_s3_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S3_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s4_sel: begin
                              m5_nxt_st[48:0] = m5_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m5_latch_cmd = m5_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m5_s4_cmd_cur = m5_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m5_s4_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S4_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s5_sel: begin
                              m5_nxt_st[48:0] = m5_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m5_latch_cmd = m5_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m5_s5_cmd_cur = m5_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m5_s5_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S5_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s6_sel: begin
                              m5_nxt_st[48:0] = m5_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m5_latch_cmd = m5_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m5_s6_cmd_cur = m5_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m5_s6_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S6_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s7_sel: begin
                              m5_nxt_st[48:0] = S_S7_DATA;
                              m5_s7_cmd_cur = 1'b1;
                             end
             m5_s7_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S7_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s8_sel: begin
                              m5_nxt_st[48:0] = m5_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m5_latch_cmd = m5_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m5_s8_cmd_cur = m5_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m5_s8_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S8_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s9_sel: begin
                              m5_nxt_st[48:0] = m5_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m5_latch_cmd = m5_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m5_s9_cmd_cur = m5_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m5_s9_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S9_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s10_sel: begin
                              m5_nxt_st[48:0] = m5_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m5_latch_cmd = m5_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m5_s10_cmd_cur = m5_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m5_s10_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S10_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s11_sel: begin
                              m5_nxt_st[48:0] = m5_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m5_latch_cmd = m5_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m5_s11_cmd_cur = m5_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m5_s11_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S11_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             default: begin
                             m5_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m5_nxt_st[48:0] = S_S7_DATA;
end
  S_S8_CMD: begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = s8_hready ? 1'b1 : 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       m5_nxt_st[48:0] = s8_hready  ? S_S8_DATA : S_S8_CMD;
  end
  S_S8_DATA:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b1;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       if(s8_hready)
         begin
           case(1'b1)
             m5_s0_sel: begin
                              m5_nxt_st[48:0] = m5_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m5_latch_cmd = m5_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m5_s0_cmd_cur = m5_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m5_s0_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S0_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s1_sel: begin
                              m5_nxt_st[48:0] = m5_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m5_latch_cmd = m5_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m5_s1_cmd_cur = m5_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m5_s1_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S1_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s2_sel: begin
                              m5_nxt_st[48:0] = m5_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m5_latch_cmd = m5_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m5_s2_cmd_cur = m5_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m5_s2_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S2_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s3_sel: begin
                              m5_nxt_st[48:0] = m5_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m5_latch_cmd = m5_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m5_s3_cmd_cur = m5_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m5_s3_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S3_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s4_sel: begin
                              m5_nxt_st[48:0] = m5_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m5_latch_cmd = m5_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m5_s4_cmd_cur = m5_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m5_s4_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S4_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s5_sel: begin
                              m5_nxt_st[48:0] = m5_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m5_latch_cmd = m5_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m5_s5_cmd_cur = m5_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m5_s5_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S5_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s6_sel: begin
                              m5_nxt_st[48:0] = m5_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m5_latch_cmd = m5_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m5_s6_cmd_cur = m5_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m5_s6_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S6_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s7_sel: begin
                              m5_nxt_st[48:0] = m5_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m5_latch_cmd = m5_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m5_s7_cmd_cur = m5_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m5_s7_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S7_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s8_sel: begin
                              m5_nxt_st[48:0] = S_S8_DATA;
                              m5_s8_cmd_cur = 1'b1;
                             end
             m5_s8_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S8_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s9_sel: begin
                              m5_nxt_st[48:0] = m5_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m5_latch_cmd = m5_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m5_s9_cmd_cur = m5_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m5_s9_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S9_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s10_sel: begin
                              m5_nxt_st[48:0] = m5_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m5_latch_cmd = m5_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m5_s10_cmd_cur = m5_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m5_s10_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S10_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s11_sel: begin
                              m5_nxt_st[48:0] = m5_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m5_latch_cmd = m5_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m5_s11_cmd_cur = m5_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m5_s11_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S11_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             default: begin
                             m5_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m5_nxt_st[48:0] = S_S8_DATA;
end
  S_S9_CMD: begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = s9_hready ? 1'b1 : 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       m5_nxt_st[48:0] = s9_hready  ? S_S9_DATA : S_S9_CMD;
  end
  S_S9_DATA:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b1;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       if(s9_hready)
         begin
           case(1'b1)
             m5_s0_sel: begin
                              m5_nxt_st[48:0] = m5_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m5_latch_cmd = m5_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m5_s0_cmd_cur = m5_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m5_s0_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S0_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s1_sel: begin
                              m5_nxt_st[48:0] = m5_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m5_latch_cmd = m5_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m5_s1_cmd_cur = m5_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m5_s1_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S1_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s2_sel: begin
                              m5_nxt_st[48:0] = m5_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m5_latch_cmd = m5_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m5_s2_cmd_cur = m5_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m5_s2_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S2_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s3_sel: begin
                              m5_nxt_st[48:0] = m5_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m5_latch_cmd = m5_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m5_s3_cmd_cur = m5_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m5_s3_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S3_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s4_sel: begin
                              m5_nxt_st[48:0] = m5_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m5_latch_cmd = m5_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m5_s4_cmd_cur = m5_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m5_s4_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S4_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s5_sel: begin
                              m5_nxt_st[48:0] = m5_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m5_latch_cmd = m5_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m5_s5_cmd_cur = m5_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m5_s5_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S5_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s6_sel: begin
                              m5_nxt_st[48:0] = m5_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m5_latch_cmd = m5_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m5_s6_cmd_cur = m5_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m5_s6_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S6_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s7_sel: begin
                              m5_nxt_st[48:0] = m5_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m5_latch_cmd = m5_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m5_s7_cmd_cur = m5_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m5_s7_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S7_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s8_sel: begin
                              m5_nxt_st[48:0] = m5_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m5_latch_cmd = m5_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m5_s8_cmd_cur = m5_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m5_s8_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S8_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s9_sel: begin
                              m5_nxt_st[48:0] = S_S9_DATA;
                              m5_s9_cmd_cur = 1'b1;
                             end
             m5_s9_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S9_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s10_sel: begin
                              m5_nxt_st[48:0] = m5_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m5_latch_cmd = m5_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m5_s10_cmd_cur = m5_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m5_s10_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S10_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s11_sel: begin
                              m5_nxt_st[48:0] = m5_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m5_latch_cmd = m5_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m5_s11_cmd_cur = m5_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m5_s11_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S11_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             default: begin
                             m5_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m5_nxt_st[48:0] = S_S9_DATA;
end
  S_S10_CMD: begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = s10_hready ? 1'b1 : 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       m5_nxt_st[48:0] = s10_hready  ? S_S10_DATA : S_S10_CMD;
  end
  S_S10_DATA:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b1;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       if(s10_hready)
         begin
           case(1'b1)
             m5_s0_sel: begin
                              m5_nxt_st[48:0] = m5_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m5_latch_cmd = m5_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m5_s0_cmd_cur = m5_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m5_s0_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S0_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s1_sel: begin
                              m5_nxt_st[48:0] = m5_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m5_latch_cmd = m5_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m5_s1_cmd_cur = m5_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m5_s1_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S1_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s2_sel: begin
                              m5_nxt_st[48:0] = m5_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m5_latch_cmd = m5_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m5_s2_cmd_cur = m5_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m5_s2_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S2_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s3_sel: begin
                              m5_nxt_st[48:0] = m5_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m5_latch_cmd = m5_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m5_s3_cmd_cur = m5_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m5_s3_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S3_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s4_sel: begin
                              m5_nxt_st[48:0] = m5_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m5_latch_cmd = m5_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m5_s4_cmd_cur = m5_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m5_s4_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S4_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s5_sel: begin
                              m5_nxt_st[48:0] = m5_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m5_latch_cmd = m5_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m5_s5_cmd_cur = m5_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m5_s5_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S5_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s6_sel: begin
                              m5_nxt_st[48:0] = m5_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m5_latch_cmd = m5_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m5_s6_cmd_cur = m5_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m5_s6_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S6_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s7_sel: begin
                              m5_nxt_st[48:0] = m5_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m5_latch_cmd = m5_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m5_s7_cmd_cur = m5_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m5_s7_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S7_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s8_sel: begin
                              m5_nxt_st[48:0] = m5_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m5_latch_cmd = m5_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m5_s8_cmd_cur = m5_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m5_s8_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S8_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s9_sel: begin
                              m5_nxt_st[48:0] = m5_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m5_latch_cmd = m5_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m5_s9_cmd_cur = m5_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m5_s9_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S9_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s10_sel: begin
                              m5_nxt_st[48:0] = S_S10_DATA;
                              m5_s10_cmd_cur = 1'b1;
                             end
             m5_s10_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S10_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s11_sel: begin
                              m5_nxt_st[48:0] = m5_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m5_latch_cmd = m5_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m5_s11_cmd_cur = m5_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m5_s11_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S11_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             default: begin
                             m5_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m5_nxt_st[48:0] = S_S10_DATA;
end
  S_S11_CMD: begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = s11_hready ? 1'b1 : 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b0;
       m5_nxt_st[48:0] = s11_hready  ? S_S11_DATA : S_S11_CMD;
  end
  S_S11_DATA:begin
       m5_latch_cmd = 1'b0;
       m5_s0_cmd_last = 1'b0;
       m5_s0_cmd_cur = 1'b0;
       m5_s0_data = 1'b0;
       m5_s1_cmd_last = 1'b0;
       m5_s1_cmd_cur = 1'b0;
       m5_s1_data = 1'b0;
       m5_s2_cmd_last = 1'b0;
       m5_s2_cmd_cur = 1'b0;
       m5_s2_data = 1'b0;
       m5_s3_cmd_last = 1'b0;
       m5_s3_cmd_cur = 1'b0;
       m5_s3_data = 1'b0;
       m5_s4_cmd_last = 1'b0;
       m5_s4_cmd_cur = 1'b0;
       m5_s4_data = 1'b0;
       m5_s5_cmd_last = 1'b0;
       m5_s5_cmd_cur = 1'b0;
       m5_s5_data = 1'b0;
       m5_s6_cmd_last = 1'b0;
       m5_s6_cmd_cur = 1'b0;
       m5_s6_data = 1'b0;
       m5_s7_cmd_last = 1'b0;
       m5_s7_cmd_cur = 1'b0;
       m5_s7_data = 1'b0;
       m5_s8_cmd_last = 1'b0;
       m5_s8_cmd_cur = 1'b0;
       m5_s8_data = 1'b0;
       m5_s9_cmd_last = 1'b0;
       m5_s9_cmd_cur = 1'b0;
       m5_s9_data = 1'b0;
       m5_s10_cmd_last = 1'b0;
       m5_s10_cmd_cur = 1'b0;
       m5_s10_data = 1'b0;
       m5_s11_cmd_last = 1'b0;
       m5_s11_cmd_cur = 1'b0;
       m5_s11_data = 1'b1;
       if(s11_hready)
         begin
           case(1'b1)
             m5_s0_sel: begin
                              m5_nxt_st[48:0] = m5_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m5_latch_cmd = m5_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m5_s0_cmd_cur = m5_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m5_s0_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S0_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s1_sel: begin
                              m5_nxt_st[48:0] = m5_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m5_latch_cmd = m5_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m5_s1_cmd_cur = m5_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m5_s1_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S1_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s2_sel: begin
                              m5_nxt_st[48:0] = m5_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m5_latch_cmd = m5_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m5_s2_cmd_cur = m5_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m5_s2_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S2_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s3_sel: begin
                              m5_nxt_st[48:0] = m5_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m5_latch_cmd = m5_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m5_s3_cmd_cur = m5_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m5_s3_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S3_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s4_sel: begin
                              m5_nxt_st[48:0] = m5_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m5_latch_cmd = m5_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m5_s4_cmd_cur = m5_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m5_s4_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S4_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s5_sel: begin
                              m5_nxt_st[48:0] = m5_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m5_latch_cmd = m5_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m5_s5_cmd_cur = m5_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m5_s5_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S5_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s6_sel: begin
                              m5_nxt_st[48:0] = m5_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m5_latch_cmd = m5_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m5_s6_cmd_cur = m5_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m5_s6_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S6_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s7_sel: begin
                              m5_nxt_st[48:0] = m5_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m5_latch_cmd = m5_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m5_s7_cmd_cur = m5_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m5_s7_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S7_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s8_sel: begin
                              m5_nxt_st[48:0] = m5_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m5_latch_cmd = m5_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m5_s8_cmd_cur = m5_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m5_s8_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S8_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s9_sel: begin
                              m5_nxt_st[48:0] = m5_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m5_latch_cmd = m5_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m5_s9_cmd_cur = m5_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m5_s9_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S9_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s10_sel: begin
                              m5_nxt_st[48:0] = m5_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m5_latch_cmd = m5_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m5_s10_cmd_cur = m5_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m5_s10_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S10_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             m5_s11_sel: begin
                              m5_nxt_st[48:0] = S_S11_DATA;
                              m5_s11_cmd_cur = 1'b1;
                             end
             m5_s11_wt_sel: begin
                                 m5_nxt_st[48:0] = S_S11_GNT;
                                 m5_latch_cmd = 1'b1;
                               end
             default: begin
                             m5_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m5_nxt_st[48:0] = S_S11_DATA;
end
  default: begin
             m5_latch_cmd = 1'b0;
             m5_s0_cmd_last = 1'b0;
             m5_s0_cmd_cur = 1'b0;
             m5_s0_data = 1'b0;
             m5_s1_cmd_last = 1'b0;
             m5_s1_cmd_cur = 1'b0;
             m5_s1_data = 1'b0;
             m5_s2_cmd_last = 1'b0;
             m5_s2_cmd_cur = 1'b0;
             m5_s2_data = 1'b0;
             m5_s3_cmd_last = 1'b0;
             m5_s3_cmd_cur = 1'b0;
             m5_s3_data = 1'b0;
             m5_s4_cmd_last = 1'b0;
             m5_s4_cmd_cur = 1'b0;
             m5_s4_data = 1'b0;
             m5_s5_cmd_last = 1'b0;
             m5_s5_cmd_cur = 1'b0;
             m5_s5_data = 1'b0;
             m5_s6_cmd_last = 1'b0;
             m5_s6_cmd_cur = 1'b0;
             m5_s6_data = 1'b0;
             m5_s7_cmd_last = 1'b0;
             m5_s7_cmd_cur = 1'b0;
             m5_s7_data = 1'b0;
             m5_s8_cmd_last = 1'b0;
             m5_s8_cmd_cur = 1'b0;
             m5_s8_data = 1'b0;
             m5_s9_cmd_last = 1'b0;
             m5_s9_cmd_cur = 1'b0;
             m5_s9_data = 1'b0;
             m5_s10_cmd_last = 1'b0;
             m5_s10_cmd_cur = 1'b0;
             m5_s10_data = 1'b0;
             m5_s11_cmd_last = 1'b0;
             m5_s11_cmd_cur = 1'b0;
             m5_s11_data = 1'b0;
             m5_nxt_st[48:0] = S_IDLE;
  end
endcase
end
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
       m6_cur_st[48:0] <= S_IDLE;
    else
       m6_cur_st[48:0] <= m6_nxt_st[48:0];
  end
always @ (*)
begin
case(m6_cur_st[48:0])
  S_IDLE:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       case(1'b1)
         m6_s0_sel: begin
                          m6_nxt_st[48:0] = m6_s0_hld ? S_S0_WAIT : (s0_hready ? S_S0_DATA : S_S0_CMD);
                          m6_latch_cmd = m6_s0_hld ? 1'b1 : (s0_hready ? 1'b0 : 1'b1);
                          m6_s0_cmd_cur = m6_s0_hld ? 1'b0 : (s0_hready ? 1'b1 : 1'b0);
                        end
         m6_s0_wt_sel: begin
                             m6_nxt_st[48:0] = S_S0_GNT;
                             m6_latch_cmd = 1'b1;
                           end
         m6_s1_sel: begin
                          m6_nxt_st[48:0] = m6_s1_hld ? S_S1_WAIT : (s1_hready ? S_S1_DATA : S_S1_CMD);
                          m6_latch_cmd = m6_s1_hld ? 1'b1 : (s1_hready ? 1'b0 : 1'b1);
                          m6_s1_cmd_cur = m6_s1_hld ? 1'b0 : (s1_hready ? 1'b1 : 1'b0);
                        end
         m6_s1_wt_sel: begin
                             m6_nxt_st[48:0] = S_S1_GNT;
                             m6_latch_cmd = 1'b1;
                           end
         m6_s2_sel: begin
                          m6_nxt_st[48:0] = m6_s2_hld ? S_S2_WAIT : (s2_hready ? S_S2_DATA : S_S2_CMD);
                          m6_latch_cmd = m6_s2_hld ? 1'b1 : (s2_hready ? 1'b0 : 1'b1);
                          m6_s2_cmd_cur = m6_s2_hld ? 1'b0 : (s2_hready ? 1'b1 : 1'b0);
                        end
         m6_s2_wt_sel: begin
                             m6_nxt_st[48:0] = S_S2_GNT;
                             m6_latch_cmd = 1'b1;
                           end
         m6_s3_sel: begin
                          m6_nxt_st[48:0] = m6_s3_hld ? S_S3_WAIT : (s3_hready ? S_S3_DATA : S_S3_CMD);
                          m6_latch_cmd = m6_s3_hld ? 1'b1 : (s3_hready ? 1'b0 : 1'b1);
                          m6_s3_cmd_cur = m6_s3_hld ? 1'b0 : (s3_hready ? 1'b1 : 1'b0);
                        end
         m6_s3_wt_sel: begin
                             m6_nxt_st[48:0] = S_S3_GNT;
                             m6_latch_cmd = 1'b1;
                           end
         m6_s4_sel: begin
                          m6_nxt_st[48:0] = m6_s4_hld ? S_S4_WAIT : (s4_hready ? S_S4_DATA : S_S4_CMD);
                          m6_latch_cmd = m6_s4_hld ? 1'b1 : (s4_hready ? 1'b0 : 1'b1);
                          m6_s4_cmd_cur = m6_s4_hld ? 1'b0 : (s4_hready ? 1'b1 : 1'b0);
                        end
         m6_s4_wt_sel: begin
                             m6_nxt_st[48:0] = S_S4_GNT;
                             m6_latch_cmd = 1'b1;
                           end
         m6_s5_sel: begin
                          m6_nxt_st[48:0] = m6_s5_hld ? S_S5_WAIT : (s5_hready ? S_S5_DATA : S_S5_CMD);
                          m6_latch_cmd = m6_s5_hld ? 1'b1 : (s5_hready ? 1'b0 : 1'b1);
                          m6_s5_cmd_cur = m6_s5_hld ? 1'b0 : (s5_hready ? 1'b1 : 1'b0);
                        end
         m6_s5_wt_sel: begin
                             m6_nxt_st[48:0] = S_S5_GNT;
                             m6_latch_cmd = 1'b1;
                           end
         m6_s6_sel: begin
                          m6_nxt_st[48:0] = m6_s6_hld ? S_S6_WAIT : (s6_hready ? S_S6_DATA : S_S6_CMD);
                          m6_latch_cmd = m6_s6_hld ? 1'b1 : (s6_hready ? 1'b0 : 1'b1);
                          m6_s6_cmd_cur = m6_s6_hld ? 1'b0 : (s6_hready ? 1'b1 : 1'b0);
                        end
         m6_s6_wt_sel: begin
                             m6_nxt_st[48:0] = S_S6_GNT;
                             m6_latch_cmd = 1'b1;
                           end
         m6_s7_sel: begin
                          m6_nxt_st[48:0] = m6_s7_hld ? S_S7_WAIT : (s7_hready ? S_S7_DATA : S_S7_CMD);
                          m6_latch_cmd = m6_s7_hld ? 1'b1 : (s7_hready ? 1'b0 : 1'b1);
                          m6_s7_cmd_cur = m6_s7_hld ? 1'b0 : (s7_hready ? 1'b1 : 1'b0);
                        end
         m6_s7_wt_sel: begin
                             m6_nxt_st[48:0] = S_S7_GNT;
                             m6_latch_cmd = 1'b1;
                           end
         m6_s8_sel: begin
                          m6_nxt_st[48:0] = m6_s8_hld ? S_S8_WAIT : (s8_hready ? S_S8_DATA : S_S8_CMD);
                          m6_latch_cmd = m6_s8_hld ? 1'b1 : (s8_hready ? 1'b0 : 1'b1);
                          m6_s8_cmd_cur = m6_s8_hld ? 1'b0 : (s8_hready ? 1'b1 : 1'b0);
                        end
         m6_s8_wt_sel: begin
                             m6_nxt_st[48:0] = S_S8_GNT;
                             m6_latch_cmd = 1'b1;
                           end
         m6_s9_sel: begin
                          m6_nxt_st[48:0] = m6_s9_hld ? S_S9_WAIT : (s9_hready ? S_S9_DATA : S_S9_CMD);
                          m6_latch_cmd = m6_s9_hld ? 1'b1 : (s9_hready ? 1'b0 : 1'b1);
                          m6_s9_cmd_cur = m6_s9_hld ? 1'b0 : (s9_hready ? 1'b1 : 1'b0);
                        end
         m6_s9_wt_sel: begin
                             m6_nxt_st[48:0] = S_S9_GNT;
                             m6_latch_cmd = 1'b1;
                           end
         m6_s10_sel: begin
                          m6_nxt_st[48:0] = m6_s10_hld ? S_S10_WAIT : (s10_hready ? S_S10_DATA : S_S10_CMD);
                          m6_latch_cmd = m6_s10_hld ? 1'b1 : (s10_hready ? 1'b0 : 1'b1);
                          m6_s10_cmd_cur = m6_s10_hld ? 1'b0 : (s10_hready ? 1'b1 : 1'b0);
                        end
         m6_s10_wt_sel: begin
                             m6_nxt_st[48:0] = S_S10_GNT;
                             m6_latch_cmd = 1'b1;
                           end
         m6_s11_sel: begin
                          m6_nxt_st[48:0] = m6_s11_hld ? S_S11_WAIT : (s11_hready ? S_S11_DATA : S_S11_CMD);
                          m6_latch_cmd = m6_s11_hld ? 1'b1 : (s11_hready ? 1'b0 : 1'b1);
                          m6_s11_cmd_cur = m6_s11_hld ? 1'b0 : (s11_hready ? 1'b1 : 1'b0);
                        end
         m6_s11_wt_sel: begin
                             m6_nxt_st[48:0] = S_S11_GNT;
                             m6_latch_cmd = 1'b1;
                           end
         default: begin
                          m6_nxt_st[48:0] = S_IDLE;
                  end
       endcase
  end
  S_S0_GNT:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       case(1'b1)
         m6_s0_sel: begin
                          m6_nxt_st[48:0] = m6_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                          m6_s0_cmd_last = m6_s0_hld ? 1'b0 : (s0_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m6_nxt_st[48:0] = S_S0_GNT;
                  end
       endcase
  end
  S_S1_GNT:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       case(1'b1)
         m6_s1_sel: begin
                          m6_nxt_st[48:0] = m6_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                          m6_s1_cmd_last = m6_s1_hld ? 1'b0 : (s1_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m6_nxt_st[48:0] = S_S1_GNT;
                  end
       endcase
  end
  S_S2_GNT:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       case(1'b1)
         m6_s2_sel: begin
                          m6_nxt_st[48:0] = m6_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                          m6_s2_cmd_last = m6_s2_hld ? 1'b0 : (s2_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m6_nxt_st[48:0] = S_S2_GNT;
                  end
       endcase
  end
  S_S3_GNT:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       case(1'b1)
         m6_s3_sel: begin
                          m6_nxt_st[48:0] = m6_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                          m6_s3_cmd_last = m6_s3_hld ? 1'b0 : (s3_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m6_nxt_st[48:0] = S_S3_GNT;
                  end
       endcase
  end
  S_S4_GNT:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       case(1'b1)
         m6_s4_sel: begin
                          m6_nxt_st[48:0] = m6_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                          m6_s4_cmd_last = m6_s4_hld ? 1'b0 : (s4_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m6_nxt_st[48:0] = S_S4_GNT;
                  end
       endcase
  end
  S_S5_GNT:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       case(1'b1)
         m6_s5_sel: begin
                          m6_nxt_st[48:0] = m6_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                          m6_s5_cmd_last = m6_s5_hld ? 1'b0 : (s5_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m6_nxt_st[48:0] = S_S5_GNT;
                  end
       endcase
  end
  S_S6_GNT:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       case(1'b1)
         m6_s6_sel: begin
                          m6_nxt_st[48:0] = m6_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                          m6_s6_cmd_last = m6_s6_hld ? 1'b0 : (s6_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m6_nxt_st[48:0] = S_S6_GNT;
                  end
       endcase
  end
  S_S7_GNT:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       case(1'b1)
         m6_s7_sel: begin
                          m6_nxt_st[48:0] = m6_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                          m6_s7_cmd_last = m6_s7_hld ? 1'b0 : (s7_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m6_nxt_st[48:0] = S_S7_GNT;
                  end
       endcase
  end
  S_S8_GNT:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       case(1'b1)
         m6_s8_sel: begin
                          m6_nxt_st[48:0] = m6_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                          m6_s8_cmd_last = m6_s8_hld ? 1'b0 : (s8_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m6_nxt_st[48:0] = S_S8_GNT;
                  end
       endcase
  end
  S_S9_GNT:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       case(1'b1)
         m6_s9_sel: begin
                          m6_nxt_st[48:0] = m6_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                          m6_s9_cmd_last = m6_s9_hld ? 1'b0 : (s9_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m6_nxt_st[48:0] = S_S9_GNT;
                  end
       endcase
  end
  S_S10_GNT:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       case(1'b1)
         m6_s10_sel: begin
                          m6_nxt_st[48:0] = m6_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                          m6_s10_cmd_last = m6_s10_hld ? 1'b0 : (s10_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m6_nxt_st[48:0] = S_S10_GNT;
                  end
       endcase
  end
  S_S11_GNT:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       case(1'b1)
         m6_s11_sel: begin
                          m6_nxt_st[48:0] = m6_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                          m6_s11_cmd_last = m6_s11_hld ? 1'b0 : (s11_hready ? 1'b1 : 1'b0);
                        end
         default: begin
                          m6_nxt_st[48:0] = S_S11_GNT;
                  end
       endcase
  end
  S_S0_WAIT:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       case(1'b1)
         ~m6_s0_hld: begin
                          m6_nxt_st[48:0] = m6_s0_wt_sel ? S_S0_GNT : s0_hready ? S_S0_DATA : S_S0_CMD;
                          m6_s0_cmd_last = m6_s0_wt_sel ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m6_nxt_st[48:0] = S_S0_WAIT;
                  end
       endcase
  end
  S_S1_WAIT:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       case(1'b1)
         ~m6_s1_hld: begin
                          m6_nxt_st[48:0] = m6_s1_wt_sel ? S_S1_GNT : s1_hready ? S_S1_DATA : S_S1_CMD;
                          m6_s1_cmd_last = m6_s1_wt_sel ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m6_nxt_st[48:0] = S_S1_WAIT;
                  end
       endcase
  end
  S_S2_WAIT:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       case(1'b1)
         ~m6_s2_hld: begin
                          m6_nxt_st[48:0] = m6_s2_wt_sel ? S_S2_GNT : s2_hready ? S_S2_DATA : S_S2_CMD;
                          m6_s2_cmd_last = m6_s2_wt_sel ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m6_nxt_st[48:0] = S_S2_WAIT;
                  end
       endcase
  end
  S_S3_WAIT:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       case(1'b1)
         ~m6_s3_hld: begin
                          m6_nxt_st[48:0] = m6_s3_wt_sel ? S_S3_GNT : s3_hready ? S_S3_DATA : S_S3_CMD;
                          m6_s3_cmd_last = m6_s3_wt_sel ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m6_nxt_st[48:0] = S_S3_WAIT;
                  end
       endcase
  end
  S_S4_WAIT:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       case(1'b1)
         ~m6_s4_hld: begin
                          m6_nxt_st[48:0] = m6_s4_wt_sel ? S_S4_GNT : s4_hready ? S_S4_DATA : S_S4_CMD;
                          m6_s4_cmd_last = m6_s4_wt_sel ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m6_nxt_st[48:0] = S_S4_WAIT;
                  end
       endcase
  end
  S_S5_WAIT:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       case(1'b1)
         ~m6_s5_hld: begin
                          m6_nxt_st[48:0] = m6_s5_wt_sel ? S_S5_GNT : s5_hready ? S_S5_DATA : S_S5_CMD;
                          m6_s5_cmd_last = m6_s5_wt_sel ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m6_nxt_st[48:0] = S_S5_WAIT;
                  end
       endcase
  end
  S_S6_WAIT:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       case(1'b1)
         ~m6_s6_hld: begin
                          m6_nxt_st[48:0] = m6_s6_wt_sel ? S_S6_GNT : s6_hready ? S_S6_DATA : S_S6_CMD;
                          m6_s6_cmd_last = m6_s6_wt_sel ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m6_nxt_st[48:0] = S_S6_WAIT;
                  end
       endcase
  end
  S_S7_WAIT:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       case(1'b1)
         ~m6_s7_hld: begin
                          m6_nxt_st[48:0] = m6_s7_wt_sel ? S_S7_GNT : s7_hready ? S_S7_DATA : S_S7_CMD;
                          m6_s7_cmd_last = m6_s7_wt_sel ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m6_nxt_st[48:0] = S_S7_WAIT;
                  end
       endcase
  end
  S_S8_WAIT:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       case(1'b1)
         ~m6_s8_hld: begin
                          m6_nxt_st[48:0] = m6_s8_wt_sel ? S_S8_GNT : s8_hready ? S_S8_DATA : S_S8_CMD;
                          m6_s8_cmd_last = m6_s8_wt_sel ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m6_nxt_st[48:0] = S_S8_WAIT;
                  end
       endcase
  end
  S_S9_WAIT:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       case(1'b1)
         ~m6_s9_hld: begin
                          m6_nxt_st[48:0] = m6_s9_wt_sel ? S_S9_GNT : s9_hready ? S_S9_DATA : S_S9_CMD;
                          m6_s9_cmd_last = m6_s9_wt_sel ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m6_nxt_st[48:0] = S_S9_WAIT;
                  end
       endcase
  end
  S_S10_WAIT:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       case(1'b1)
         ~m6_s10_hld: begin
                          m6_nxt_st[48:0] = m6_s10_wt_sel ? S_S10_GNT : s10_hready ? S_S10_DATA : S_S10_CMD;
                          m6_s10_cmd_last = m6_s10_wt_sel ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m6_nxt_st[48:0] = S_S10_WAIT;
                  end
       endcase
  end
  S_S11_WAIT:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       case(1'b1)
         ~m6_s11_hld: begin
                          m6_nxt_st[48:0] = m6_s11_wt_sel ? S_S11_GNT : s11_hready ? S_S11_DATA : S_S11_CMD;
                          m6_s11_cmd_last = m6_s11_wt_sel ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                        end
         default: begin
                          m6_nxt_st[48:0] = S_S11_WAIT;
                  end
       endcase
  end
  S_S0_CMD: begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = s0_hready ? 1'b1 : 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       m6_nxt_st[48:0] = s0_hready  ? S_S0_DATA : S_S0_CMD;
  end
  S_S0_DATA:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b1;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       if(s0_hready)
         begin
           case(1'b1)
             m6_s0_sel: begin
                              m6_nxt_st[48:0] = S_S0_DATA;
                              m6_s0_cmd_cur = 1'b1;
                             end
             m6_s0_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S0_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s1_sel: begin
                              m6_nxt_st[48:0] = m6_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m6_latch_cmd = m6_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m6_s1_cmd_cur = m6_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m6_s1_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S1_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s2_sel: begin
                              m6_nxt_st[48:0] = m6_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m6_latch_cmd = m6_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m6_s2_cmd_cur = m6_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m6_s2_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S2_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s3_sel: begin
                              m6_nxt_st[48:0] = m6_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m6_latch_cmd = m6_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m6_s3_cmd_cur = m6_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m6_s3_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S3_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s4_sel: begin
                              m6_nxt_st[48:0] = m6_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m6_latch_cmd = m6_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m6_s4_cmd_cur = m6_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m6_s4_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S4_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s5_sel: begin
                              m6_nxt_st[48:0] = m6_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m6_latch_cmd = m6_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m6_s5_cmd_cur = m6_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m6_s5_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S5_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s6_sel: begin
                              m6_nxt_st[48:0] = m6_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m6_latch_cmd = m6_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m6_s6_cmd_cur = m6_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m6_s6_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S6_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s7_sel: begin
                              m6_nxt_st[48:0] = m6_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m6_latch_cmd = m6_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m6_s7_cmd_cur = m6_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m6_s7_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S7_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s8_sel: begin
                              m6_nxt_st[48:0] = m6_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m6_latch_cmd = m6_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m6_s8_cmd_cur = m6_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m6_s8_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S8_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s9_sel: begin
                              m6_nxt_st[48:0] = m6_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m6_latch_cmd = m6_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m6_s9_cmd_cur = m6_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m6_s9_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S9_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s10_sel: begin
                              m6_nxt_st[48:0] = m6_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m6_latch_cmd = m6_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m6_s10_cmd_cur = m6_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m6_s10_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S10_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s11_sel: begin
                              m6_nxt_st[48:0] = m6_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m6_latch_cmd = m6_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m6_s11_cmd_cur = m6_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m6_s11_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S11_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             default: begin
                             m6_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m6_nxt_st[48:0] = S_S0_DATA;
end
  S_S1_CMD: begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = s1_hready ? 1'b1 : 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       m6_nxt_st[48:0] = s1_hready  ? S_S1_DATA : S_S1_CMD;
  end
  S_S1_DATA:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b1;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       if(s1_hready)
         begin
           case(1'b1)
             m6_s0_sel: begin
                              m6_nxt_st[48:0] = m6_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m6_latch_cmd = m6_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m6_s0_cmd_cur = m6_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m6_s0_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S0_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s1_sel: begin
                              m6_nxt_st[48:0] = S_S1_DATA;
                              m6_s1_cmd_cur = 1'b1;
                             end
             m6_s1_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S1_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s2_sel: begin
                              m6_nxt_st[48:0] = m6_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m6_latch_cmd = m6_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m6_s2_cmd_cur = m6_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m6_s2_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S2_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s3_sel: begin
                              m6_nxt_st[48:0] = m6_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m6_latch_cmd = m6_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m6_s3_cmd_cur = m6_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m6_s3_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S3_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s4_sel: begin
                              m6_nxt_st[48:0] = m6_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m6_latch_cmd = m6_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m6_s4_cmd_cur = m6_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m6_s4_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S4_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s5_sel: begin
                              m6_nxt_st[48:0] = m6_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m6_latch_cmd = m6_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m6_s5_cmd_cur = m6_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m6_s5_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S5_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s6_sel: begin
                              m6_nxt_st[48:0] = m6_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m6_latch_cmd = m6_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m6_s6_cmd_cur = m6_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m6_s6_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S6_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s7_sel: begin
                              m6_nxt_st[48:0] = m6_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m6_latch_cmd = m6_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m6_s7_cmd_cur = m6_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m6_s7_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S7_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s8_sel: begin
                              m6_nxt_st[48:0] = m6_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m6_latch_cmd = m6_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m6_s8_cmd_cur = m6_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m6_s8_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S8_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s9_sel: begin
                              m6_nxt_st[48:0] = m6_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m6_latch_cmd = m6_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m6_s9_cmd_cur = m6_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m6_s9_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S9_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s10_sel: begin
                              m6_nxt_st[48:0] = m6_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m6_latch_cmd = m6_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m6_s10_cmd_cur = m6_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m6_s10_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S10_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s11_sel: begin
                              m6_nxt_st[48:0] = m6_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m6_latch_cmd = m6_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m6_s11_cmd_cur = m6_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m6_s11_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S11_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             default: begin
                             m6_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m6_nxt_st[48:0] = S_S1_DATA;
end
  S_S2_CMD: begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = s2_hready ? 1'b1 : 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       m6_nxt_st[48:0] = s2_hready  ? S_S2_DATA : S_S2_CMD;
  end
  S_S2_DATA:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b1;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       if(s2_hready)
         begin
           case(1'b1)
             m6_s0_sel: begin
                              m6_nxt_st[48:0] = m6_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m6_latch_cmd = m6_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m6_s0_cmd_cur = m6_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m6_s0_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S0_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s1_sel: begin
                              m6_nxt_st[48:0] = m6_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m6_latch_cmd = m6_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m6_s1_cmd_cur = m6_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m6_s1_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S1_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s2_sel: begin
                              m6_nxt_st[48:0] = S_S2_DATA;
                              m6_s2_cmd_cur = 1'b1;
                             end
             m6_s2_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S2_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s3_sel: begin
                              m6_nxt_st[48:0] = m6_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m6_latch_cmd = m6_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m6_s3_cmd_cur = m6_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m6_s3_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S3_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s4_sel: begin
                              m6_nxt_st[48:0] = m6_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m6_latch_cmd = m6_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m6_s4_cmd_cur = m6_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m6_s4_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S4_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s5_sel: begin
                              m6_nxt_st[48:0] = m6_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m6_latch_cmd = m6_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m6_s5_cmd_cur = m6_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m6_s5_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S5_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s6_sel: begin
                              m6_nxt_st[48:0] = m6_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m6_latch_cmd = m6_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m6_s6_cmd_cur = m6_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m6_s6_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S6_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s7_sel: begin
                              m6_nxt_st[48:0] = m6_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m6_latch_cmd = m6_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m6_s7_cmd_cur = m6_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m6_s7_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S7_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s8_sel: begin
                              m6_nxt_st[48:0] = m6_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m6_latch_cmd = m6_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m6_s8_cmd_cur = m6_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m6_s8_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S8_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s9_sel: begin
                              m6_nxt_st[48:0] = m6_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m6_latch_cmd = m6_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m6_s9_cmd_cur = m6_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m6_s9_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S9_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s10_sel: begin
                              m6_nxt_st[48:0] = m6_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m6_latch_cmd = m6_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m6_s10_cmd_cur = m6_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m6_s10_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S10_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s11_sel: begin
                              m6_nxt_st[48:0] = m6_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m6_latch_cmd = m6_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m6_s11_cmd_cur = m6_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m6_s11_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S11_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             default: begin
                             m6_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m6_nxt_st[48:0] = S_S2_DATA;
end
  S_S3_CMD: begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = s3_hready ? 1'b1 : 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       m6_nxt_st[48:0] = s3_hready  ? S_S3_DATA : S_S3_CMD;
  end
  S_S3_DATA:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b1;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       if(s3_hready)
         begin
           case(1'b1)
             m6_s0_sel: begin
                              m6_nxt_st[48:0] = m6_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m6_latch_cmd = m6_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m6_s0_cmd_cur = m6_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m6_s0_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S0_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s1_sel: begin
                              m6_nxt_st[48:0] = m6_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m6_latch_cmd = m6_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m6_s1_cmd_cur = m6_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m6_s1_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S1_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s2_sel: begin
                              m6_nxt_st[48:0] = m6_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m6_latch_cmd = m6_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m6_s2_cmd_cur = m6_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m6_s2_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S2_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s3_sel: begin
                              m6_nxt_st[48:0] = S_S3_DATA;
                              m6_s3_cmd_cur = 1'b1;
                             end
             m6_s3_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S3_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s4_sel: begin
                              m6_nxt_st[48:0] = m6_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m6_latch_cmd = m6_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m6_s4_cmd_cur = m6_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m6_s4_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S4_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s5_sel: begin
                              m6_nxt_st[48:0] = m6_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m6_latch_cmd = m6_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m6_s5_cmd_cur = m6_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m6_s5_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S5_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s6_sel: begin
                              m6_nxt_st[48:0] = m6_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m6_latch_cmd = m6_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m6_s6_cmd_cur = m6_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m6_s6_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S6_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s7_sel: begin
                              m6_nxt_st[48:0] = m6_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m6_latch_cmd = m6_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m6_s7_cmd_cur = m6_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m6_s7_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S7_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s8_sel: begin
                              m6_nxt_st[48:0] = m6_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m6_latch_cmd = m6_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m6_s8_cmd_cur = m6_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m6_s8_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S8_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s9_sel: begin
                              m6_nxt_st[48:0] = m6_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m6_latch_cmd = m6_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m6_s9_cmd_cur = m6_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m6_s9_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S9_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s10_sel: begin
                              m6_nxt_st[48:0] = m6_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m6_latch_cmd = m6_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m6_s10_cmd_cur = m6_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m6_s10_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S10_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s11_sel: begin
                              m6_nxt_st[48:0] = m6_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m6_latch_cmd = m6_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m6_s11_cmd_cur = m6_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m6_s11_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S11_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             default: begin
                             m6_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m6_nxt_st[48:0] = S_S3_DATA;
end
  S_S4_CMD: begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = s4_hready ? 1'b1 : 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       m6_nxt_st[48:0] = s4_hready  ? S_S4_DATA : S_S4_CMD;
  end
  S_S4_DATA:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b1;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       if(s4_hready)
         begin
           case(1'b1)
             m6_s0_sel: begin
                              m6_nxt_st[48:0] = m6_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m6_latch_cmd = m6_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m6_s0_cmd_cur = m6_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m6_s0_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S0_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s1_sel: begin
                              m6_nxt_st[48:0] = m6_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m6_latch_cmd = m6_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m6_s1_cmd_cur = m6_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m6_s1_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S1_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s2_sel: begin
                              m6_nxt_st[48:0] = m6_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m6_latch_cmd = m6_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m6_s2_cmd_cur = m6_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m6_s2_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S2_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s3_sel: begin
                              m6_nxt_st[48:0] = m6_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m6_latch_cmd = m6_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m6_s3_cmd_cur = m6_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m6_s3_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S3_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s4_sel: begin
                              m6_nxt_st[48:0] = S_S4_DATA;
                              m6_s4_cmd_cur = 1'b1;
                             end
             m6_s4_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S4_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s5_sel: begin
                              m6_nxt_st[48:0] = m6_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m6_latch_cmd = m6_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m6_s5_cmd_cur = m6_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m6_s5_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S5_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s6_sel: begin
                              m6_nxt_st[48:0] = m6_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m6_latch_cmd = m6_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m6_s6_cmd_cur = m6_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m6_s6_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S6_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s7_sel: begin
                              m6_nxt_st[48:0] = m6_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m6_latch_cmd = m6_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m6_s7_cmd_cur = m6_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m6_s7_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S7_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s8_sel: begin
                              m6_nxt_st[48:0] = m6_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m6_latch_cmd = m6_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m6_s8_cmd_cur = m6_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m6_s8_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S8_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s9_sel: begin
                              m6_nxt_st[48:0] = m6_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m6_latch_cmd = m6_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m6_s9_cmd_cur = m6_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m6_s9_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S9_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s10_sel: begin
                              m6_nxt_st[48:0] = m6_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m6_latch_cmd = m6_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m6_s10_cmd_cur = m6_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m6_s10_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S10_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s11_sel: begin
                              m6_nxt_st[48:0] = m6_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m6_latch_cmd = m6_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m6_s11_cmd_cur = m6_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m6_s11_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S11_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             default: begin
                             m6_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m6_nxt_st[48:0] = S_S4_DATA;
end
  S_S5_CMD: begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = s5_hready ? 1'b1 : 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       m6_nxt_st[48:0] = s5_hready  ? S_S5_DATA : S_S5_CMD;
  end
  S_S5_DATA:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b1;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       if(s5_hready)
         begin
           case(1'b1)
             m6_s0_sel: begin
                              m6_nxt_st[48:0] = m6_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m6_latch_cmd = m6_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m6_s0_cmd_cur = m6_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m6_s0_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S0_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s1_sel: begin
                              m6_nxt_st[48:0] = m6_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m6_latch_cmd = m6_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m6_s1_cmd_cur = m6_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m6_s1_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S1_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s2_sel: begin
                              m6_nxt_st[48:0] = m6_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m6_latch_cmd = m6_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m6_s2_cmd_cur = m6_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m6_s2_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S2_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s3_sel: begin
                              m6_nxt_st[48:0] = m6_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m6_latch_cmd = m6_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m6_s3_cmd_cur = m6_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m6_s3_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S3_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s4_sel: begin
                              m6_nxt_st[48:0] = m6_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m6_latch_cmd = m6_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m6_s4_cmd_cur = m6_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m6_s4_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S4_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s5_sel: begin
                              m6_nxt_st[48:0] = S_S5_DATA;
                              m6_s5_cmd_cur = 1'b1;
                             end
             m6_s5_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S5_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s6_sel: begin
                              m6_nxt_st[48:0] = m6_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m6_latch_cmd = m6_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m6_s6_cmd_cur = m6_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m6_s6_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S6_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s7_sel: begin
                              m6_nxt_st[48:0] = m6_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m6_latch_cmd = m6_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m6_s7_cmd_cur = m6_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m6_s7_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S7_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s8_sel: begin
                              m6_nxt_st[48:0] = m6_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m6_latch_cmd = m6_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m6_s8_cmd_cur = m6_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m6_s8_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S8_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s9_sel: begin
                              m6_nxt_st[48:0] = m6_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m6_latch_cmd = m6_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m6_s9_cmd_cur = m6_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m6_s9_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S9_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s10_sel: begin
                              m6_nxt_st[48:0] = m6_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m6_latch_cmd = m6_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m6_s10_cmd_cur = m6_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m6_s10_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S10_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s11_sel: begin
                              m6_nxt_st[48:0] = m6_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m6_latch_cmd = m6_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m6_s11_cmd_cur = m6_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m6_s11_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S11_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             default: begin
                             m6_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m6_nxt_st[48:0] = S_S5_DATA;
end
  S_S6_CMD: begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = s6_hready ? 1'b1 : 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       m6_nxt_st[48:0] = s6_hready  ? S_S6_DATA : S_S6_CMD;
  end
  S_S6_DATA:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b1;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       if(s6_hready)
         begin
           case(1'b1)
             m6_s0_sel: begin
                              m6_nxt_st[48:0] = m6_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m6_latch_cmd = m6_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m6_s0_cmd_cur = m6_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m6_s0_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S0_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s1_sel: begin
                              m6_nxt_st[48:0] = m6_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m6_latch_cmd = m6_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m6_s1_cmd_cur = m6_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m6_s1_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S1_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s2_sel: begin
                              m6_nxt_st[48:0] = m6_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m6_latch_cmd = m6_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m6_s2_cmd_cur = m6_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m6_s2_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S2_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s3_sel: begin
                              m6_nxt_st[48:0] = m6_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m6_latch_cmd = m6_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m6_s3_cmd_cur = m6_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m6_s3_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S3_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s4_sel: begin
                              m6_nxt_st[48:0] = m6_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m6_latch_cmd = m6_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m6_s4_cmd_cur = m6_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m6_s4_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S4_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s5_sel: begin
                              m6_nxt_st[48:0] = m6_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m6_latch_cmd = m6_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m6_s5_cmd_cur = m6_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m6_s5_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S5_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s6_sel: begin
                              m6_nxt_st[48:0] = S_S6_DATA;
                              m6_s6_cmd_cur = 1'b1;
                             end
             m6_s6_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S6_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s7_sel: begin
                              m6_nxt_st[48:0] = m6_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m6_latch_cmd = m6_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m6_s7_cmd_cur = m6_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m6_s7_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S7_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s8_sel: begin
                              m6_nxt_st[48:0] = m6_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m6_latch_cmd = m6_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m6_s8_cmd_cur = m6_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m6_s8_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S8_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s9_sel: begin
                              m6_nxt_st[48:0] = m6_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m6_latch_cmd = m6_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m6_s9_cmd_cur = m6_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m6_s9_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S9_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s10_sel: begin
                              m6_nxt_st[48:0] = m6_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m6_latch_cmd = m6_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m6_s10_cmd_cur = m6_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m6_s10_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S10_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s11_sel: begin
                              m6_nxt_st[48:0] = m6_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m6_latch_cmd = m6_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m6_s11_cmd_cur = m6_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m6_s11_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S11_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             default: begin
                             m6_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m6_nxt_st[48:0] = S_S6_DATA;
end
  S_S7_CMD: begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = s7_hready ? 1'b1 : 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       m6_nxt_st[48:0] = s7_hready  ? S_S7_DATA : S_S7_CMD;
  end
  S_S7_DATA:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b1;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       if(s7_hready)
         begin
           case(1'b1)
             m6_s0_sel: begin
                              m6_nxt_st[48:0] = m6_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m6_latch_cmd = m6_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m6_s0_cmd_cur = m6_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m6_s0_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S0_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s1_sel: begin
                              m6_nxt_st[48:0] = m6_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m6_latch_cmd = m6_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m6_s1_cmd_cur = m6_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m6_s1_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S1_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s2_sel: begin
                              m6_nxt_st[48:0] = m6_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m6_latch_cmd = m6_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m6_s2_cmd_cur = m6_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m6_s2_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S2_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s3_sel: begin
                              m6_nxt_st[48:0] = m6_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m6_latch_cmd = m6_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m6_s3_cmd_cur = m6_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m6_s3_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S3_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s4_sel: begin
                              m6_nxt_st[48:0] = m6_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m6_latch_cmd = m6_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m6_s4_cmd_cur = m6_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m6_s4_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S4_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s5_sel: begin
                              m6_nxt_st[48:0] = m6_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m6_latch_cmd = m6_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m6_s5_cmd_cur = m6_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m6_s5_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S5_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s6_sel: begin
                              m6_nxt_st[48:0] = m6_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m6_latch_cmd = m6_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m6_s6_cmd_cur = m6_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m6_s6_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S6_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s7_sel: begin
                              m6_nxt_st[48:0] = S_S7_DATA;
                              m6_s7_cmd_cur = 1'b1;
                             end
             m6_s7_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S7_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s8_sel: begin
                              m6_nxt_st[48:0] = m6_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m6_latch_cmd = m6_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m6_s8_cmd_cur = m6_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m6_s8_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S8_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s9_sel: begin
                              m6_nxt_st[48:0] = m6_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m6_latch_cmd = m6_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m6_s9_cmd_cur = m6_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m6_s9_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S9_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s10_sel: begin
                              m6_nxt_st[48:0] = m6_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m6_latch_cmd = m6_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m6_s10_cmd_cur = m6_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m6_s10_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S10_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s11_sel: begin
                              m6_nxt_st[48:0] = m6_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m6_latch_cmd = m6_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m6_s11_cmd_cur = m6_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m6_s11_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S11_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             default: begin
                             m6_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m6_nxt_st[48:0] = S_S7_DATA;
end
  S_S8_CMD: begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = s8_hready ? 1'b1 : 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       m6_nxt_st[48:0] = s8_hready  ? S_S8_DATA : S_S8_CMD;
  end
  S_S8_DATA:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b1;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       if(s8_hready)
         begin
           case(1'b1)
             m6_s0_sel: begin
                              m6_nxt_st[48:0] = m6_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m6_latch_cmd = m6_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m6_s0_cmd_cur = m6_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m6_s0_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S0_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s1_sel: begin
                              m6_nxt_st[48:0] = m6_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m6_latch_cmd = m6_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m6_s1_cmd_cur = m6_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m6_s1_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S1_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s2_sel: begin
                              m6_nxt_st[48:0] = m6_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m6_latch_cmd = m6_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m6_s2_cmd_cur = m6_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m6_s2_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S2_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s3_sel: begin
                              m6_nxt_st[48:0] = m6_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m6_latch_cmd = m6_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m6_s3_cmd_cur = m6_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m6_s3_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S3_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s4_sel: begin
                              m6_nxt_st[48:0] = m6_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m6_latch_cmd = m6_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m6_s4_cmd_cur = m6_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m6_s4_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S4_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s5_sel: begin
                              m6_nxt_st[48:0] = m6_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m6_latch_cmd = m6_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m6_s5_cmd_cur = m6_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m6_s5_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S5_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s6_sel: begin
                              m6_nxt_st[48:0] = m6_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m6_latch_cmd = m6_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m6_s6_cmd_cur = m6_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m6_s6_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S6_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s7_sel: begin
                              m6_nxt_st[48:0] = m6_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m6_latch_cmd = m6_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m6_s7_cmd_cur = m6_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m6_s7_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S7_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s8_sel: begin
                              m6_nxt_st[48:0] = S_S8_DATA;
                              m6_s8_cmd_cur = 1'b1;
                             end
             m6_s8_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S8_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s9_sel: begin
                              m6_nxt_st[48:0] = m6_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m6_latch_cmd = m6_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m6_s9_cmd_cur = m6_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m6_s9_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S9_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s10_sel: begin
                              m6_nxt_st[48:0] = m6_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m6_latch_cmd = m6_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m6_s10_cmd_cur = m6_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m6_s10_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S10_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s11_sel: begin
                              m6_nxt_st[48:0] = m6_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m6_latch_cmd = m6_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m6_s11_cmd_cur = m6_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m6_s11_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S11_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             default: begin
                             m6_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m6_nxt_st[48:0] = S_S8_DATA;
end
  S_S9_CMD: begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = s9_hready ? 1'b1 : 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       m6_nxt_st[48:0] = s9_hready  ? S_S9_DATA : S_S9_CMD;
  end
  S_S9_DATA:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b1;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       if(s9_hready)
         begin
           case(1'b1)
             m6_s0_sel: begin
                              m6_nxt_st[48:0] = m6_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m6_latch_cmd = m6_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m6_s0_cmd_cur = m6_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m6_s0_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S0_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s1_sel: begin
                              m6_nxt_st[48:0] = m6_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m6_latch_cmd = m6_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m6_s1_cmd_cur = m6_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m6_s1_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S1_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s2_sel: begin
                              m6_nxt_st[48:0] = m6_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m6_latch_cmd = m6_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m6_s2_cmd_cur = m6_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m6_s2_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S2_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s3_sel: begin
                              m6_nxt_st[48:0] = m6_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m6_latch_cmd = m6_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m6_s3_cmd_cur = m6_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m6_s3_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S3_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s4_sel: begin
                              m6_nxt_st[48:0] = m6_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m6_latch_cmd = m6_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m6_s4_cmd_cur = m6_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m6_s4_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S4_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s5_sel: begin
                              m6_nxt_st[48:0] = m6_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m6_latch_cmd = m6_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m6_s5_cmd_cur = m6_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m6_s5_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S5_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s6_sel: begin
                              m6_nxt_st[48:0] = m6_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m6_latch_cmd = m6_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m6_s6_cmd_cur = m6_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m6_s6_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S6_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s7_sel: begin
                              m6_nxt_st[48:0] = m6_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m6_latch_cmd = m6_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m6_s7_cmd_cur = m6_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m6_s7_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S7_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s8_sel: begin
                              m6_nxt_st[48:0] = m6_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m6_latch_cmd = m6_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m6_s8_cmd_cur = m6_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m6_s8_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S8_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s9_sel: begin
                              m6_nxt_st[48:0] = S_S9_DATA;
                              m6_s9_cmd_cur = 1'b1;
                             end
             m6_s9_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S9_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s10_sel: begin
                              m6_nxt_st[48:0] = m6_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m6_latch_cmd = m6_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m6_s10_cmd_cur = m6_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m6_s10_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S10_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s11_sel: begin
                              m6_nxt_st[48:0] = m6_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m6_latch_cmd = m6_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m6_s11_cmd_cur = m6_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m6_s11_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S11_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             default: begin
                             m6_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m6_nxt_st[48:0] = S_S9_DATA;
end
  S_S10_CMD: begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = s10_hready ? 1'b1 : 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       m6_nxt_st[48:0] = s10_hready  ? S_S10_DATA : S_S10_CMD;
  end
  S_S10_DATA:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b1;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       if(s10_hready)
         begin
           case(1'b1)
             m6_s0_sel: begin
                              m6_nxt_st[48:0] = m6_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m6_latch_cmd = m6_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m6_s0_cmd_cur = m6_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m6_s0_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S0_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s1_sel: begin
                              m6_nxt_st[48:0] = m6_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m6_latch_cmd = m6_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m6_s1_cmd_cur = m6_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m6_s1_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S1_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s2_sel: begin
                              m6_nxt_st[48:0] = m6_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m6_latch_cmd = m6_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m6_s2_cmd_cur = m6_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m6_s2_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S2_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s3_sel: begin
                              m6_nxt_st[48:0] = m6_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m6_latch_cmd = m6_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m6_s3_cmd_cur = m6_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m6_s3_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S3_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s4_sel: begin
                              m6_nxt_st[48:0] = m6_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m6_latch_cmd = m6_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m6_s4_cmd_cur = m6_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m6_s4_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S4_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s5_sel: begin
                              m6_nxt_st[48:0] = m6_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m6_latch_cmd = m6_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m6_s5_cmd_cur = m6_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m6_s5_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S5_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s6_sel: begin
                              m6_nxt_st[48:0] = m6_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m6_latch_cmd = m6_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m6_s6_cmd_cur = m6_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m6_s6_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S6_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s7_sel: begin
                              m6_nxt_st[48:0] = m6_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m6_latch_cmd = m6_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m6_s7_cmd_cur = m6_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m6_s7_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S7_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s8_sel: begin
                              m6_nxt_st[48:0] = m6_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m6_latch_cmd = m6_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m6_s8_cmd_cur = m6_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m6_s8_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S8_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s9_sel: begin
                              m6_nxt_st[48:0] = m6_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m6_latch_cmd = m6_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m6_s9_cmd_cur = m6_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m6_s9_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S9_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s10_sel: begin
                              m6_nxt_st[48:0] = S_S10_DATA;
                              m6_s10_cmd_cur = 1'b1;
                             end
             m6_s10_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S10_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s11_sel: begin
                              m6_nxt_st[48:0] = m6_s11_hld ? S_S11_WAIT : s11_hready ? S_S11_DATA : S_S11_CMD;
                              m6_latch_cmd = m6_s11_hld ? 1'b1 : s11_hready ? 1'b0 : 1'b1;
                              m6_s11_cmd_cur = m6_s11_hld ? 1'b0 : s11_hready ? 1'b1 : 1'b0;
                            end
             m6_s11_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S11_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             default: begin
                             m6_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m6_nxt_st[48:0] = S_S10_DATA;
end
  S_S11_CMD: begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = s11_hready ? 1'b1 : 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b0;
       m6_nxt_st[48:0] = s11_hready  ? S_S11_DATA : S_S11_CMD;
  end
  S_S11_DATA:begin
       m6_latch_cmd = 1'b0;
       m6_s0_cmd_last = 1'b0;
       m6_s0_cmd_cur = 1'b0;
       m6_s0_data = 1'b0;
       m6_s1_cmd_last = 1'b0;
       m6_s1_cmd_cur = 1'b0;
       m6_s1_data = 1'b0;
       m6_s2_cmd_last = 1'b0;
       m6_s2_cmd_cur = 1'b0;
       m6_s2_data = 1'b0;
       m6_s3_cmd_last = 1'b0;
       m6_s3_cmd_cur = 1'b0;
       m6_s3_data = 1'b0;
       m6_s4_cmd_last = 1'b0;
       m6_s4_cmd_cur = 1'b0;
       m6_s4_data = 1'b0;
       m6_s5_cmd_last = 1'b0;
       m6_s5_cmd_cur = 1'b0;
       m6_s5_data = 1'b0;
       m6_s6_cmd_last = 1'b0;
       m6_s6_cmd_cur = 1'b0;
       m6_s6_data = 1'b0;
       m6_s7_cmd_last = 1'b0;
       m6_s7_cmd_cur = 1'b0;
       m6_s7_data = 1'b0;
       m6_s8_cmd_last = 1'b0;
       m6_s8_cmd_cur = 1'b0;
       m6_s8_data = 1'b0;
       m6_s9_cmd_last = 1'b0;
       m6_s9_cmd_cur = 1'b0;
       m6_s9_data = 1'b0;
       m6_s10_cmd_last = 1'b0;
       m6_s10_cmd_cur = 1'b0;
       m6_s10_data = 1'b0;
       m6_s11_cmd_last = 1'b0;
       m6_s11_cmd_cur = 1'b0;
       m6_s11_data = 1'b1;
       if(s11_hready)
         begin
           case(1'b1)
             m6_s0_sel: begin
                              m6_nxt_st[48:0] = m6_s0_hld ? S_S0_WAIT : s0_hready ? S_S0_DATA : S_S0_CMD;
                              m6_latch_cmd = m6_s0_hld ? 1'b1 : s0_hready ? 1'b0 : 1'b1;
                              m6_s0_cmd_cur = m6_s0_hld ? 1'b0 : s0_hready ? 1'b1 : 1'b0;
                            end
             m6_s0_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S0_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s1_sel: begin
                              m6_nxt_st[48:0] = m6_s1_hld ? S_S1_WAIT : s1_hready ? S_S1_DATA : S_S1_CMD;
                              m6_latch_cmd = m6_s1_hld ? 1'b1 : s1_hready ? 1'b0 : 1'b1;
                              m6_s1_cmd_cur = m6_s1_hld ? 1'b0 : s1_hready ? 1'b1 : 1'b0;
                            end
             m6_s1_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S1_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s2_sel: begin
                              m6_nxt_st[48:0] = m6_s2_hld ? S_S2_WAIT : s2_hready ? S_S2_DATA : S_S2_CMD;
                              m6_latch_cmd = m6_s2_hld ? 1'b1 : s2_hready ? 1'b0 : 1'b1;
                              m6_s2_cmd_cur = m6_s2_hld ? 1'b0 : s2_hready ? 1'b1 : 1'b0;
                            end
             m6_s2_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S2_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s3_sel: begin
                              m6_nxt_st[48:0] = m6_s3_hld ? S_S3_WAIT : s3_hready ? S_S3_DATA : S_S3_CMD;
                              m6_latch_cmd = m6_s3_hld ? 1'b1 : s3_hready ? 1'b0 : 1'b1;
                              m6_s3_cmd_cur = m6_s3_hld ? 1'b0 : s3_hready ? 1'b1 : 1'b0;
                            end
             m6_s3_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S3_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s4_sel: begin
                              m6_nxt_st[48:0] = m6_s4_hld ? S_S4_WAIT : s4_hready ? S_S4_DATA : S_S4_CMD;
                              m6_latch_cmd = m6_s4_hld ? 1'b1 : s4_hready ? 1'b0 : 1'b1;
                              m6_s4_cmd_cur = m6_s4_hld ? 1'b0 : s4_hready ? 1'b1 : 1'b0;
                            end
             m6_s4_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S4_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s5_sel: begin
                              m6_nxt_st[48:0] = m6_s5_hld ? S_S5_WAIT : s5_hready ? S_S5_DATA : S_S5_CMD;
                              m6_latch_cmd = m6_s5_hld ? 1'b1 : s5_hready ? 1'b0 : 1'b1;
                              m6_s5_cmd_cur = m6_s5_hld ? 1'b0 : s5_hready ? 1'b1 : 1'b0;
                            end
             m6_s5_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S5_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s6_sel: begin
                              m6_nxt_st[48:0] = m6_s6_hld ? S_S6_WAIT : s6_hready ? S_S6_DATA : S_S6_CMD;
                              m6_latch_cmd = m6_s6_hld ? 1'b1 : s6_hready ? 1'b0 : 1'b1;
                              m6_s6_cmd_cur = m6_s6_hld ? 1'b0 : s6_hready ? 1'b1 : 1'b0;
                            end
             m6_s6_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S6_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s7_sel: begin
                              m6_nxt_st[48:0] = m6_s7_hld ? S_S7_WAIT : s7_hready ? S_S7_DATA : S_S7_CMD;
                              m6_latch_cmd = m6_s7_hld ? 1'b1 : s7_hready ? 1'b0 : 1'b1;
                              m6_s7_cmd_cur = m6_s7_hld ? 1'b0 : s7_hready ? 1'b1 : 1'b0;
                            end
             m6_s7_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S7_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s8_sel: begin
                              m6_nxt_st[48:0] = m6_s8_hld ? S_S8_WAIT : s8_hready ? S_S8_DATA : S_S8_CMD;
                              m6_latch_cmd = m6_s8_hld ? 1'b1 : s8_hready ? 1'b0 : 1'b1;
                              m6_s8_cmd_cur = m6_s8_hld ? 1'b0 : s8_hready ? 1'b1 : 1'b0;
                            end
             m6_s8_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S8_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s9_sel: begin
                              m6_nxt_st[48:0] = m6_s9_hld ? S_S9_WAIT : s9_hready ? S_S9_DATA : S_S9_CMD;
                              m6_latch_cmd = m6_s9_hld ? 1'b1 : s9_hready ? 1'b0 : 1'b1;
                              m6_s9_cmd_cur = m6_s9_hld ? 1'b0 : s9_hready ? 1'b1 : 1'b0;
                            end
             m6_s9_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S9_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s10_sel: begin
                              m6_nxt_st[48:0] = m6_s10_hld ? S_S10_WAIT : s10_hready ? S_S10_DATA : S_S10_CMD;
                              m6_latch_cmd = m6_s10_hld ? 1'b1 : s10_hready ? 1'b0 : 1'b1;
                              m6_s10_cmd_cur = m6_s10_hld ? 1'b0 : s10_hready ? 1'b1 : 1'b0;
                            end
             m6_s10_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S10_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             m6_s11_sel: begin
                              m6_nxt_st[48:0] = S_S11_DATA;
                              m6_s11_cmd_cur = 1'b1;
                             end
             m6_s11_wt_sel: begin
                                 m6_nxt_st[48:0] = S_S11_GNT;
                                 m6_latch_cmd = 1'b1;
                               end
             default: begin
                             m6_nxt_st[48:0] = S_IDLE;
                      end
           endcase
         end
       else
         m6_nxt_st[48:0] = S_S11_DATA;
end
  default: begin
             m6_latch_cmd = 1'b0;
             m6_s0_cmd_last = 1'b0;
             m6_s0_cmd_cur = 1'b0;
             m6_s0_data = 1'b0;
             m6_s1_cmd_last = 1'b0;
             m6_s1_cmd_cur = 1'b0;
             m6_s1_data = 1'b0;
             m6_s2_cmd_last = 1'b0;
             m6_s2_cmd_cur = 1'b0;
             m6_s2_data = 1'b0;
             m6_s3_cmd_last = 1'b0;
             m6_s3_cmd_cur = 1'b0;
             m6_s3_data = 1'b0;
             m6_s4_cmd_last = 1'b0;
             m6_s4_cmd_cur = 1'b0;
             m6_s4_data = 1'b0;
             m6_s5_cmd_last = 1'b0;
             m6_s5_cmd_cur = 1'b0;
             m6_s5_data = 1'b0;
             m6_s6_cmd_last = 1'b0;
             m6_s6_cmd_cur = 1'b0;
             m6_s6_data = 1'b0;
             m6_s7_cmd_last = 1'b0;
             m6_s7_cmd_cur = 1'b0;
             m6_s7_data = 1'b0;
             m6_s8_cmd_last = 1'b0;
             m6_s8_cmd_cur = 1'b0;
             m6_s8_data = 1'b0;
             m6_s9_cmd_last = 1'b0;
             m6_s9_cmd_cur = 1'b0;
             m6_s9_data = 1'b0;
             m6_s10_cmd_last = 1'b0;
             m6_s10_cmd_cur = 1'b0;
             m6_s10_data = 1'b0;
             m6_s11_cmd_last = 1'b0;
             m6_s11_cmd_cur = 1'b0;
             m6_s11_data = 1'b0;
             m6_nxt_st[48:0] = S_IDLE;
  end
endcase
end
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m0_s0_req_pend_tmp <= 1'b0;
    else if(m0_latch_cmd && m0_s0_req)
        m0_s0_req_pend_tmp <= 1'b1;
    else if((m0_cur_st[48:0] == S_S0_DATA) && s0_hready)
        m0_s0_req_pend_tmp <= 1'b0;
  end
assign m0_s0_req_pend = m0_s0_req_pend_tmp && (~((m0_cur_st[48:0] == S_S0_DATA) && s0_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m0_s1_req_pend_tmp <= 1'b0;
    else if(m0_latch_cmd && m0_s1_req)
        m0_s1_req_pend_tmp <= 1'b1;
    else if((m0_cur_st[48:0] == S_S1_DATA) && s1_hready)
        m0_s1_req_pend_tmp <= 1'b0;
  end
assign m0_s1_req_pend = m0_s1_req_pend_tmp && (~((m0_cur_st[48:0] == S_S1_DATA) && s1_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m0_s2_req_pend_tmp <= 1'b0;
    else if(m0_latch_cmd && m0_s2_req)
        m0_s2_req_pend_tmp <= 1'b1;
    else if((m0_cur_st[48:0] == S_S2_DATA) && s2_hready)
        m0_s2_req_pend_tmp <= 1'b0;
  end
assign m0_s2_req_pend = m0_s2_req_pend_tmp && (~((m0_cur_st[48:0] == S_S2_DATA) && s2_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m0_s3_req_pend_tmp <= 1'b0;
    else if(m0_latch_cmd && m0_s3_req)
        m0_s3_req_pend_tmp <= 1'b1;
    else if((m0_cur_st[48:0] == S_S3_DATA) && s3_hready)
        m0_s3_req_pend_tmp <= 1'b0;
  end
assign m0_s3_req_pend = m0_s3_req_pend_tmp && (~((m0_cur_st[48:0] == S_S3_DATA) && s3_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m0_s4_req_pend_tmp <= 1'b0;
    else if(m0_latch_cmd && m0_s4_req)
        m0_s4_req_pend_tmp <= 1'b1;
    else if((m0_cur_st[48:0] == S_S4_DATA) && s4_hready)
        m0_s4_req_pend_tmp <= 1'b0;
  end
assign m0_s4_req_pend = m0_s4_req_pend_tmp && (~((m0_cur_st[48:0] == S_S4_DATA) && s4_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m0_s5_req_pend_tmp <= 1'b0;
    else if(m0_latch_cmd && m0_s5_req)
        m0_s5_req_pend_tmp <= 1'b1;
    else if((m0_cur_st[48:0] == S_S5_DATA) && s5_hready)
        m0_s5_req_pend_tmp <= 1'b0;
  end
assign m0_s5_req_pend = m0_s5_req_pend_tmp && (~((m0_cur_st[48:0] == S_S5_DATA) && s5_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m0_s6_req_pend_tmp <= 1'b0;
    else if(m0_latch_cmd && m0_s6_req)
        m0_s6_req_pend_tmp <= 1'b1;
    else if((m0_cur_st[48:0] == S_S6_DATA) && s6_hready)
        m0_s6_req_pend_tmp <= 1'b0;
  end
assign m0_s6_req_pend = m0_s6_req_pend_tmp && (~((m0_cur_st[48:0] == S_S6_DATA) && s6_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m0_s7_req_pend_tmp <= 1'b0;
    else if(m0_latch_cmd && m0_s7_req)
        m0_s7_req_pend_tmp <= 1'b1;
    else if((m0_cur_st[48:0] == S_S7_DATA) && s7_hready)
        m0_s7_req_pend_tmp <= 1'b0;
  end
assign m0_s7_req_pend = m0_s7_req_pend_tmp && (~((m0_cur_st[48:0] == S_S7_DATA) && s7_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m0_s8_req_pend_tmp <= 1'b0;
    else if(m0_latch_cmd && m0_s8_req)
        m0_s8_req_pend_tmp <= 1'b1;
    else if((m0_cur_st[48:0] == S_S8_DATA) && s8_hready)
        m0_s8_req_pend_tmp <= 1'b0;
  end
assign m0_s8_req_pend = m0_s8_req_pend_tmp && (~((m0_cur_st[48:0] == S_S8_DATA) && s8_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m0_s9_req_pend_tmp <= 1'b0;
    else if(m0_latch_cmd && m0_s9_req)
        m0_s9_req_pend_tmp <= 1'b1;
    else if((m0_cur_st[48:0] == S_S9_DATA) && s9_hready)
        m0_s9_req_pend_tmp <= 1'b0;
  end
assign m0_s9_req_pend = m0_s9_req_pend_tmp && (~((m0_cur_st[48:0] == S_S9_DATA) && s9_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m0_s10_req_pend_tmp <= 1'b0;
    else if(m0_latch_cmd && m0_s10_req)
        m0_s10_req_pend_tmp <= 1'b1;
    else if((m0_cur_st[48:0] == S_S10_DATA) && s10_hready)
        m0_s10_req_pend_tmp <= 1'b0;
  end
assign m0_s10_req_pend = m0_s10_req_pend_tmp && (~((m0_cur_st[48:0] == S_S10_DATA) && s10_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m0_s11_req_pend_tmp <= 1'b0;
    else if(m0_latch_cmd && m0_s11_req)
        m0_s11_req_pend_tmp <= 1'b1;
    else if((m0_cur_st[48:0] == S_S11_DATA) && s11_hready)
        m0_s11_req_pend_tmp <= 1'b0;
  end
assign m0_s11_req_pend = m0_s11_req_pend_tmp && (~((m0_cur_st[48:0] == S_S11_DATA) && s11_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m1_s0_req_pend_tmp <= 1'b0;
    else if(m1_latch_cmd && m1_s0_req)
        m1_s0_req_pend_tmp <= 1'b1;
    else if((m1_cur_st[48:0] == S_S0_DATA) && s0_hready)
        m1_s0_req_pend_tmp <= 1'b0;
  end
assign m1_s0_req_pend = m1_s0_req_pend_tmp && (~((m1_cur_st[48:0] == S_S0_DATA) && s0_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m1_s1_req_pend_tmp <= 1'b0;
    else if(m1_latch_cmd && m1_s1_req)
        m1_s1_req_pend_tmp <= 1'b1;
    else if((m1_cur_st[48:0] == S_S1_DATA) && s1_hready)
        m1_s1_req_pend_tmp <= 1'b0;
  end
assign m1_s1_req_pend = m1_s1_req_pend_tmp && (~((m1_cur_st[48:0] == S_S1_DATA) && s1_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m1_s2_req_pend_tmp <= 1'b0;
    else if(m1_latch_cmd && m1_s2_req)
        m1_s2_req_pend_tmp <= 1'b1;
    else if((m1_cur_st[48:0] == S_S2_DATA) && s2_hready)
        m1_s2_req_pend_tmp <= 1'b0;
  end
assign m1_s2_req_pend = m1_s2_req_pend_tmp && (~((m1_cur_st[48:0] == S_S2_DATA) && s2_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m1_s3_req_pend_tmp <= 1'b0;
    else if(m1_latch_cmd && m1_s3_req)
        m1_s3_req_pend_tmp <= 1'b1;
    else if((m1_cur_st[48:0] == S_S3_DATA) && s3_hready)
        m1_s3_req_pend_tmp <= 1'b0;
  end
assign m1_s3_req_pend = m1_s3_req_pend_tmp && (~((m1_cur_st[48:0] == S_S3_DATA) && s3_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m1_s4_req_pend_tmp <= 1'b0;
    else if(m1_latch_cmd && m1_s4_req)
        m1_s4_req_pend_tmp <= 1'b1;
    else if((m1_cur_st[48:0] == S_S4_DATA) && s4_hready)
        m1_s4_req_pend_tmp <= 1'b0;
  end
assign m1_s4_req_pend = m1_s4_req_pend_tmp && (~((m1_cur_st[48:0] == S_S4_DATA) && s4_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m1_s5_req_pend_tmp <= 1'b0;
    else if(m1_latch_cmd && m1_s5_req)
        m1_s5_req_pend_tmp <= 1'b1;
    else if((m1_cur_st[48:0] == S_S5_DATA) && s5_hready)
        m1_s5_req_pend_tmp <= 1'b0;
  end
assign m1_s5_req_pend = m1_s5_req_pend_tmp && (~((m1_cur_st[48:0] == S_S5_DATA) && s5_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m1_s6_req_pend_tmp <= 1'b0;
    else if(m1_latch_cmd && m1_s6_req)
        m1_s6_req_pend_tmp <= 1'b1;
    else if((m1_cur_st[48:0] == S_S6_DATA) && s6_hready)
        m1_s6_req_pend_tmp <= 1'b0;
  end
assign m1_s6_req_pend = m1_s6_req_pend_tmp && (~((m1_cur_st[48:0] == S_S6_DATA) && s6_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m1_s7_req_pend_tmp <= 1'b0;
    else if(m1_latch_cmd && m1_s7_req)
        m1_s7_req_pend_tmp <= 1'b1;
    else if((m1_cur_st[48:0] == S_S7_DATA) && s7_hready)
        m1_s7_req_pend_tmp <= 1'b0;
  end
assign m1_s7_req_pend = m1_s7_req_pend_tmp && (~((m1_cur_st[48:0] == S_S7_DATA) && s7_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m1_s8_req_pend_tmp <= 1'b0;
    else if(m1_latch_cmd && m1_s8_req)
        m1_s8_req_pend_tmp <= 1'b1;
    else if((m1_cur_st[48:0] == S_S8_DATA) && s8_hready)
        m1_s8_req_pend_tmp <= 1'b0;
  end
assign m1_s8_req_pend = m1_s8_req_pend_tmp && (~((m1_cur_st[48:0] == S_S8_DATA) && s8_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m1_s9_req_pend_tmp <= 1'b0;
    else if(m1_latch_cmd && m1_s9_req)
        m1_s9_req_pend_tmp <= 1'b1;
    else if((m1_cur_st[48:0] == S_S9_DATA) && s9_hready)
        m1_s9_req_pend_tmp <= 1'b0;
  end
assign m1_s9_req_pend = m1_s9_req_pend_tmp && (~((m1_cur_st[48:0] == S_S9_DATA) && s9_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m1_s10_req_pend_tmp <= 1'b0;
    else if(m1_latch_cmd && m1_s10_req)
        m1_s10_req_pend_tmp <= 1'b1;
    else if((m1_cur_st[48:0] == S_S10_DATA) && s10_hready)
        m1_s10_req_pend_tmp <= 1'b0;
  end
assign m1_s10_req_pend = m1_s10_req_pend_tmp && (~((m1_cur_st[48:0] == S_S10_DATA) && s10_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m1_s11_req_pend_tmp <= 1'b0;
    else if(m1_latch_cmd && m1_s11_req)
        m1_s11_req_pend_tmp <= 1'b1;
    else if((m1_cur_st[48:0] == S_S11_DATA) && s11_hready)
        m1_s11_req_pend_tmp <= 1'b0;
  end
assign m1_s11_req_pend = m1_s11_req_pend_tmp && (~((m1_cur_st[48:0] == S_S11_DATA) && s11_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m2_s0_req_pend_tmp <= 1'b0;
    else if(m2_latch_cmd && m2_s0_req)
        m2_s0_req_pend_tmp <= 1'b1;
    else if((m2_cur_st[48:0] == S_S0_DATA) && s0_hready)
        m2_s0_req_pend_tmp <= 1'b0;
  end
assign m2_s0_req_pend = m2_s0_req_pend_tmp && (~((m2_cur_st[48:0] == S_S0_DATA) && s0_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m2_s1_req_pend_tmp <= 1'b0;
    else if(m2_latch_cmd && m2_s1_req)
        m2_s1_req_pend_tmp <= 1'b1;
    else if((m2_cur_st[48:0] == S_S1_DATA) && s1_hready)
        m2_s1_req_pend_tmp <= 1'b0;
  end
assign m2_s1_req_pend = m2_s1_req_pend_tmp && (~((m2_cur_st[48:0] == S_S1_DATA) && s1_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m2_s2_req_pend_tmp <= 1'b0;
    else if(m2_latch_cmd && m2_s2_req)
        m2_s2_req_pend_tmp <= 1'b1;
    else if((m2_cur_st[48:0] == S_S2_DATA) && s2_hready)
        m2_s2_req_pend_tmp <= 1'b0;
  end
assign m2_s2_req_pend = m2_s2_req_pend_tmp && (~((m2_cur_st[48:0] == S_S2_DATA) && s2_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m2_s3_req_pend_tmp <= 1'b0;
    else if(m2_latch_cmd && m2_s3_req)
        m2_s3_req_pend_tmp <= 1'b1;
    else if((m2_cur_st[48:0] == S_S3_DATA) && s3_hready)
        m2_s3_req_pend_tmp <= 1'b0;
  end
assign m2_s3_req_pend = m2_s3_req_pend_tmp && (~((m2_cur_st[48:0] == S_S3_DATA) && s3_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m2_s4_req_pend_tmp <= 1'b0;
    else if(m2_latch_cmd && m2_s4_req)
        m2_s4_req_pend_tmp <= 1'b1;
    else if((m2_cur_st[48:0] == S_S4_DATA) && s4_hready)
        m2_s4_req_pend_tmp <= 1'b0;
  end
assign m2_s4_req_pend = m2_s4_req_pend_tmp && (~((m2_cur_st[48:0] == S_S4_DATA) && s4_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m2_s5_req_pend_tmp <= 1'b0;
    else if(m2_latch_cmd && m2_s5_req)
        m2_s5_req_pend_tmp <= 1'b1;
    else if((m2_cur_st[48:0] == S_S5_DATA) && s5_hready)
        m2_s5_req_pend_tmp <= 1'b0;
  end
assign m2_s5_req_pend = m2_s5_req_pend_tmp && (~((m2_cur_st[48:0] == S_S5_DATA) && s5_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m2_s6_req_pend_tmp <= 1'b0;
    else if(m2_latch_cmd && m2_s6_req)
        m2_s6_req_pend_tmp <= 1'b1;
    else if((m2_cur_st[48:0] == S_S6_DATA) && s6_hready)
        m2_s6_req_pend_tmp <= 1'b0;
  end
assign m2_s6_req_pend = m2_s6_req_pend_tmp && (~((m2_cur_st[48:0] == S_S6_DATA) && s6_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m2_s7_req_pend_tmp <= 1'b0;
    else if(m2_latch_cmd && m2_s7_req)
        m2_s7_req_pend_tmp <= 1'b1;
    else if((m2_cur_st[48:0] == S_S7_DATA) && s7_hready)
        m2_s7_req_pend_tmp <= 1'b0;
  end
assign m2_s7_req_pend = m2_s7_req_pend_tmp && (~((m2_cur_st[48:0] == S_S7_DATA) && s7_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m2_s8_req_pend_tmp <= 1'b0;
    else if(m2_latch_cmd && m2_s8_req)
        m2_s8_req_pend_tmp <= 1'b1;
    else if((m2_cur_st[48:0] == S_S8_DATA) && s8_hready)
        m2_s8_req_pend_tmp <= 1'b0;
  end
assign m2_s8_req_pend = m2_s8_req_pend_tmp && (~((m2_cur_st[48:0] == S_S8_DATA) && s8_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m2_s9_req_pend_tmp <= 1'b0;
    else if(m2_latch_cmd && m2_s9_req)
        m2_s9_req_pend_tmp <= 1'b1;
    else if((m2_cur_st[48:0] == S_S9_DATA) && s9_hready)
        m2_s9_req_pend_tmp <= 1'b0;
  end
assign m2_s9_req_pend = m2_s9_req_pend_tmp && (~((m2_cur_st[48:0] == S_S9_DATA) && s9_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m2_s10_req_pend_tmp <= 1'b0;
    else if(m2_latch_cmd && m2_s10_req)
        m2_s10_req_pend_tmp <= 1'b1;
    else if((m2_cur_st[48:0] == S_S10_DATA) && s10_hready)
        m2_s10_req_pend_tmp <= 1'b0;
  end
assign m2_s10_req_pend = m2_s10_req_pend_tmp && (~((m2_cur_st[48:0] == S_S10_DATA) && s10_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m2_s11_req_pend_tmp <= 1'b0;
    else if(m2_latch_cmd && m2_s11_req)
        m2_s11_req_pend_tmp <= 1'b1;
    else if((m2_cur_st[48:0] == S_S11_DATA) && s11_hready)
        m2_s11_req_pend_tmp <= 1'b0;
  end
assign m2_s11_req_pend = m2_s11_req_pend_tmp && (~((m2_cur_st[48:0] == S_S11_DATA) && s11_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m3_s0_req_pend_tmp <= 1'b0;
    else if(m3_latch_cmd && m3_s0_req)
        m3_s0_req_pend_tmp <= 1'b1;
    else if((m3_cur_st[48:0] == S_S0_DATA) && s0_hready)
        m3_s0_req_pend_tmp <= 1'b0;
  end
assign m3_s0_req_pend = m3_s0_req_pend_tmp && (~((m3_cur_st[48:0] == S_S0_DATA) && s0_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m3_s1_req_pend_tmp <= 1'b0;
    else if(m3_latch_cmd && m3_s1_req)
        m3_s1_req_pend_tmp <= 1'b1;
    else if((m3_cur_st[48:0] == S_S1_DATA) && s1_hready)
        m3_s1_req_pend_tmp <= 1'b0;
  end
assign m3_s1_req_pend = m3_s1_req_pend_tmp && (~((m3_cur_st[48:0] == S_S1_DATA) && s1_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m3_s2_req_pend_tmp <= 1'b0;
    else if(m3_latch_cmd && m3_s2_req)
        m3_s2_req_pend_tmp <= 1'b1;
    else if((m3_cur_st[48:0] == S_S2_DATA) && s2_hready)
        m3_s2_req_pend_tmp <= 1'b0;
  end
assign m3_s2_req_pend = m3_s2_req_pend_tmp && (~((m3_cur_st[48:0] == S_S2_DATA) && s2_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m3_s3_req_pend_tmp <= 1'b0;
    else if(m3_latch_cmd && m3_s3_req)
        m3_s3_req_pend_tmp <= 1'b1;
    else if((m3_cur_st[48:0] == S_S3_DATA) && s3_hready)
        m3_s3_req_pend_tmp <= 1'b0;
  end
assign m3_s3_req_pend = m3_s3_req_pend_tmp && (~((m3_cur_st[48:0] == S_S3_DATA) && s3_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m3_s4_req_pend_tmp <= 1'b0;
    else if(m3_latch_cmd && m3_s4_req)
        m3_s4_req_pend_tmp <= 1'b1;
    else if((m3_cur_st[48:0] == S_S4_DATA) && s4_hready)
        m3_s4_req_pend_tmp <= 1'b0;
  end
assign m3_s4_req_pend = m3_s4_req_pend_tmp && (~((m3_cur_st[48:0] == S_S4_DATA) && s4_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m3_s5_req_pend_tmp <= 1'b0;
    else if(m3_latch_cmd && m3_s5_req)
        m3_s5_req_pend_tmp <= 1'b1;
    else if((m3_cur_st[48:0] == S_S5_DATA) && s5_hready)
        m3_s5_req_pend_tmp <= 1'b0;
  end
assign m3_s5_req_pend = m3_s5_req_pend_tmp && (~((m3_cur_st[48:0] == S_S5_DATA) && s5_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m3_s6_req_pend_tmp <= 1'b0;
    else if(m3_latch_cmd && m3_s6_req)
        m3_s6_req_pend_tmp <= 1'b1;
    else if((m3_cur_st[48:0] == S_S6_DATA) && s6_hready)
        m3_s6_req_pend_tmp <= 1'b0;
  end
assign m3_s6_req_pend = m3_s6_req_pend_tmp && (~((m3_cur_st[48:0] == S_S6_DATA) && s6_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m3_s7_req_pend_tmp <= 1'b0;
    else if(m3_latch_cmd && m3_s7_req)
        m3_s7_req_pend_tmp <= 1'b1;
    else if((m3_cur_st[48:0] == S_S7_DATA) && s7_hready)
        m3_s7_req_pend_tmp <= 1'b0;
  end
assign m3_s7_req_pend = m3_s7_req_pend_tmp && (~((m3_cur_st[48:0] == S_S7_DATA) && s7_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m3_s8_req_pend_tmp <= 1'b0;
    else if(m3_latch_cmd && m3_s8_req)
        m3_s8_req_pend_tmp <= 1'b1;
    else if((m3_cur_st[48:0] == S_S8_DATA) && s8_hready)
        m3_s8_req_pend_tmp <= 1'b0;
  end
assign m3_s8_req_pend = m3_s8_req_pend_tmp && (~((m3_cur_st[48:0] == S_S8_DATA) && s8_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m3_s9_req_pend_tmp <= 1'b0;
    else if(m3_latch_cmd && m3_s9_req)
        m3_s9_req_pend_tmp <= 1'b1;
    else if((m3_cur_st[48:0] == S_S9_DATA) && s9_hready)
        m3_s9_req_pend_tmp <= 1'b0;
  end
assign m3_s9_req_pend = m3_s9_req_pend_tmp && (~((m3_cur_st[48:0] == S_S9_DATA) && s9_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m3_s10_req_pend_tmp <= 1'b0;
    else if(m3_latch_cmd && m3_s10_req)
        m3_s10_req_pend_tmp <= 1'b1;
    else if((m3_cur_st[48:0] == S_S10_DATA) && s10_hready)
        m3_s10_req_pend_tmp <= 1'b0;
  end
assign m3_s10_req_pend = m3_s10_req_pend_tmp && (~((m3_cur_st[48:0] == S_S10_DATA) && s10_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m3_s11_req_pend_tmp <= 1'b0;
    else if(m3_latch_cmd && m3_s11_req)
        m3_s11_req_pend_tmp <= 1'b1;
    else if((m3_cur_st[48:0] == S_S11_DATA) && s11_hready)
        m3_s11_req_pend_tmp <= 1'b0;
  end
assign m3_s11_req_pend = m3_s11_req_pend_tmp && (~((m3_cur_st[48:0] == S_S11_DATA) && s11_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m4_s0_req_pend_tmp <= 1'b0;
    else if(m4_latch_cmd && m4_s0_req)
        m4_s0_req_pend_tmp <= 1'b1;
    else if((m4_cur_st[48:0] == S_S0_DATA) && s0_hready)
        m4_s0_req_pend_tmp <= 1'b0;
  end
assign m4_s0_req_pend = m4_s0_req_pend_tmp && (~((m4_cur_st[48:0] == S_S0_DATA) && s0_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m4_s1_req_pend_tmp <= 1'b0;
    else if(m4_latch_cmd && m4_s1_req)
        m4_s1_req_pend_tmp <= 1'b1;
    else if((m4_cur_st[48:0] == S_S1_DATA) && s1_hready)
        m4_s1_req_pend_tmp <= 1'b0;
  end
assign m4_s1_req_pend = m4_s1_req_pend_tmp && (~((m4_cur_st[48:0] == S_S1_DATA) && s1_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m4_s2_req_pend_tmp <= 1'b0;
    else if(m4_latch_cmd && m4_s2_req)
        m4_s2_req_pend_tmp <= 1'b1;
    else if((m4_cur_st[48:0] == S_S2_DATA) && s2_hready)
        m4_s2_req_pend_tmp <= 1'b0;
  end
assign m4_s2_req_pend = m4_s2_req_pend_tmp && (~((m4_cur_st[48:0] == S_S2_DATA) && s2_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m4_s3_req_pend_tmp <= 1'b0;
    else if(m4_latch_cmd && m4_s3_req)
        m4_s3_req_pend_tmp <= 1'b1;
    else if((m4_cur_st[48:0] == S_S3_DATA) && s3_hready)
        m4_s3_req_pend_tmp <= 1'b0;
  end
assign m4_s3_req_pend = m4_s3_req_pend_tmp && (~((m4_cur_st[48:0] == S_S3_DATA) && s3_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m4_s4_req_pend_tmp <= 1'b0;
    else if(m4_latch_cmd && m4_s4_req)
        m4_s4_req_pend_tmp <= 1'b1;
    else if((m4_cur_st[48:0] == S_S4_DATA) && s4_hready)
        m4_s4_req_pend_tmp <= 1'b0;
  end
assign m4_s4_req_pend = m4_s4_req_pend_tmp && (~((m4_cur_st[48:0] == S_S4_DATA) && s4_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m4_s5_req_pend_tmp <= 1'b0;
    else if(m4_latch_cmd && m4_s5_req)
        m4_s5_req_pend_tmp <= 1'b1;
    else if((m4_cur_st[48:0] == S_S5_DATA) && s5_hready)
        m4_s5_req_pend_tmp <= 1'b0;
  end
assign m4_s5_req_pend = m4_s5_req_pend_tmp && (~((m4_cur_st[48:0] == S_S5_DATA) && s5_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m4_s6_req_pend_tmp <= 1'b0;
    else if(m4_latch_cmd && m4_s6_req)
        m4_s6_req_pend_tmp <= 1'b1;
    else if((m4_cur_st[48:0] == S_S6_DATA) && s6_hready)
        m4_s6_req_pend_tmp <= 1'b0;
  end
assign m4_s6_req_pend = m4_s6_req_pend_tmp && (~((m4_cur_st[48:0] == S_S6_DATA) && s6_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m4_s7_req_pend_tmp <= 1'b0;
    else if(m4_latch_cmd && m4_s7_req)
        m4_s7_req_pend_tmp <= 1'b1;
    else if((m4_cur_st[48:0] == S_S7_DATA) && s7_hready)
        m4_s7_req_pend_tmp <= 1'b0;
  end
assign m4_s7_req_pend = m4_s7_req_pend_tmp && (~((m4_cur_st[48:0] == S_S7_DATA) && s7_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m4_s8_req_pend_tmp <= 1'b0;
    else if(m4_latch_cmd && m4_s8_req)
        m4_s8_req_pend_tmp <= 1'b1;
    else if((m4_cur_st[48:0] == S_S8_DATA) && s8_hready)
        m4_s8_req_pend_tmp <= 1'b0;
  end
assign m4_s8_req_pend = m4_s8_req_pend_tmp && (~((m4_cur_st[48:0] == S_S8_DATA) && s8_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m4_s9_req_pend_tmp <= 1'b0;
    else if(m4_latch_cmd && m4_s9_req)
        m4_s9_req_pend_tmp <= 1'b1;
    else if((m4_cur_st[48:0] == S_S9_DATA) && s9_hready)
        m4_s9_req_pend_tmp <= 1'b0;
  end
assign m4_s9_req_pend = m4_s9_req_pend_tmp && (~((m4_cur_st[48:0] == S_S9_DATA) && s9_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m4_s10_req_pend_tmp <= 1'b0;
    else if(m4_latch_cmd && m4_s10_req)
        m4_s10_req_pend_tmp <= 1'b1;
    else if((m4_cur_st[48:0] == S_S10_DATA) && s10_hready)
        m4_s10_req_pend_tmp <= 1'b0;
  end
assign m4_s10_req_pend = m4_s10_req_pend_tmp && (~((m4_cur_st[48:0] == S_S10_DATA) && s10_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m4_s11_req_pend_tmp <= 1'b0;
    else if(m4_latch_cmd && m4_s11_req)
        m4_s11_req_pend_tmp <= 1'b1;
    else if((m4_cur_st[48:0] == S_S11_DATA) && s11_hready)
        m4_s11_req_pend_tmp <= 1'b0;
  end
assign m4_s11_req_pend = m4_s11_req_pend_tmp && (~((m4_cur_st[48:0] == S_S11_DATA) && s11_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m5_s0_req_pend_tmp <= 1'b0;
    else if(m5_latch_cmd && m5_s0_req)
        m5_s0_req_pend_tmp <= 1'b1;
    else if((m5_cur_st[48:0] == S_S0_DATA) && s0_hready)
        m5_s0_req_pend_tmp <= 1'b0;
  end
assign m5_s0_req_pend = m5_s0_req_pend_tmp && (~((m5_cur_st[48:0] == S_S0_DATA) && s0_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m5_s1_req_pend_tmp <= 1'b0;
    else if(m5_latch_cmd && m5_s1_req)
        m5_s1_req_pend_tmp <= 1'b1;
    else if((m5_cur_st[48:0] == S_S1_DATA) && s1_hready)
        m5_s1_req_pend_tmp <= 1'b0;
  end
assign m5_s1_req_pend = m5_s1_req_pend_tmp && (~((m5_cur_st[48:0] == S_S1_DATA) && s1_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m5_s2_req_pend_tmp <= 1'b0;
    else if(m5_latch_cmd && m5_s2_req)
        m5_s2_req_pend_tmp <= 1'b1;
    else if((m5_cur_st[48:0] == S_S2_DATA) && s2_hready)
        m5_s2_req_pend_tmp <= 1'b0;
  end
assign m5_s2_req_pend = m5_s2_req_pend_tmp && (~((m5_cur_st[48:0] == S_S2_DATA) && s2_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m5_s3_req_pend_tmp <= 1'b0;
    else if(m5_latch_cmd && m5_s3_req)
        m5_s3_req_pend_tmp <= 1'b1;
    else if((m5_cur_st[48:0] == S_S3_DATA) && s3_hready)
        m5_s3_req_pend_tmp <= 1'b0;
  end
assign m5_s3_req_pend = m5_s3_req_pend_tmp && (~((m5_cur_st[48:0] == S_S3_DATA) && s3_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m5_s4_req_pend_tmp <= 1'b0;
    else if(m5_latch_cmd && m5_s4_req)
        m5_s4_req_pend_tmp <= 1'b1;
    else if((m5_cur_st[48:0] == S_S4_DATA) && s4_hready)
        m5_s4_req_pend_tmp <= 1'b0;
  end
assign m5_s4_req_pend = m5_s4_req_pend_tmp && (~((m5_cur_st[48:0] == S_S4_DATA) && s4_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m5_s5_req_pend_tmp <= 1'b0;
    else if(m5_latch_cmd && m5_s5_req)
        m5_s5_req_pend_tmp <= 1'b1;
    else if((m5_cur_st[48:0] == S_S5_DATA) && s5_hready)
        m5_s5_req_pend_tmp <= 1'b0;
  end
assign m5_s5_req_pend = m5_s5_req_pend_tmp && (~((m5_cur_st[48:0] == S_S5_DATA) && s5_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m5_s6_req_pend_tmp <= 1'b0;
    else if(m5_latch_cmd && m5_s6_req)
        m5_s6_req_pend_tmp <= 1'b1;
    else if((m5_cur_st[48:0] == S_S6_DATA) && s6_hready)
        m5_s6_req_pend_tmp <= 1'b0;
  end
assign m5_s6_req_pend = m5_s6_req_pend_tmp && (~((m5_cur_st[48:0] == S_S6_DATA) && s6_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m5_s7_req_pend_tmp <= 1'b0;
    else if(m5_latch_cmd && m5_s7_req)
        m5_s7_req_pend_tmp <= 1'b1;
    else if((m5_cur_st[48:0] == S_S7_DATA) && s7_hready)
        m5_s7_req_pend_tmp <= 1'b0;
  end
assign m5_s7_req_pend = m5_s7_req_pend_tmp && (~((m5_cur_st[48:0] == S_S7_DATA) && s7_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m5_s8_req_pend_tmp <= 1'b0;
    else if(m5_latch_cmd && m5_s8_req)
        m5_s8_req_pend_tmp <= 1'b1;
    else if((m5_cur_st[48:0] == S_S8_DATA) && s8_hready)
        m5_s8_req_pend_tmp <= 1'b0;
  end
assign m5_s8_req_pend = m5_s8_req_pend_tmp && (~((m5_cur_st[48:0] == S_S8_DATA) && s8_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m5_s9_req_pend_tmp <= 1'b0;
    else if(m5_latch_cmd && m5_s9_req)
        m5_s9_req_pend_tmp <= 1'b1;
    else if((m5_cur_st[48:0] == S_S9_DATA) && s9_hready)
        m5_s9_req_pend_tmp <= 1'b0;
  end
assign m5_s9_req_pend = m5_s9_req_pend_tmp && (~((m5_cur_st[48:0] == S_S9_DATA) && s9_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m5_s10_req_pend_tmp <= 1'b0;
    else if(m5_latch_cmd && m5_s10_req)
        m5_s10_req_pend_tmp <= 1'b1;
    else if((m5_cur_st[48:0] == S_S10_DATA) && s10_hready)
        m5_s10_req_pend_tmp <= 1'b0;
  end
assign m5_s10_req_pend = m5_s10_req_pend_tmp && (~((m5_cur_st[48:0] == S_S10_DATA) && s10_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m5_s11_req_pend_tmp <= 1'b0;
    else if(m5_latch_cmd && m5_s11_req)
        m5_s11_req_pend_tmp <= 1'b1;
    else if((m5_cur_st[48:0] == S_S11_DATA) && s11_hready)
        m5_s11_req_pend_tmp <= 1'b0;
  end
assign m5_s11_req_pend = m5_s11_req_pend_tmp && (~((m5_cur_st[48:0] == S_S11_DATA) && s11_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m6_s0_req_pend_tmp <= 1'b0;
    else if(m6_latch_cmd && m6_s0_req)
        m6_s0_req_pend_tmp <= 1'b1;
    else if((m6_cur_st[48:0] == S_S0_DATA) && s0_hready)
        m6_s0_req_pend_tmp <= 1'b0;
  end
assign m6_s0_req_pend = m6_s0_req_pend_tmp && (~((m6_cur_st[48:0] == S_S0_DATA) && s0_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m6_s1_req_pend_tmp <= 1'b0;
    else if(m6_latch_cmd && m6_s1_req)
        m6_s1_req_pend_tmp <= 1'b1;
    else if((m6_cur_st[48:0] == S_S1_DATA) && s1_hready)
        m6_s1_req_pend_tmp <= 1'b0;
  end
assign m6_s1_req_pend = m6_s1_req_pend_tmp && (~((m6_cur_st[48:0] == S_S1_DATA) && s1_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m6_s2_req_pend_tmp <= 1'b0;
    else if(m6_latch_cmd && m6_s2_req)
        m6_s2_req_pend_tmp <= 1'b1;
    else if((m6_cur_st[48:0] == S_S2_DATA) && s2_hready)
        m6_s2_req_pend_tmp <= 1'b0;
  end
assign m6_s2_req_pend = m6_s2_req_pend_tmp && (~((m6_cur_st[48:0] == S_S2_DATA) && s2_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m6_s3_req_pend_tmp <= 1'b0;
    else if(m6_latch_cmd && m6_s3_req)
        m6_s3_req_pend_tmp <= 1'b1;
    else if((m6_cur_st[48:0] == S_S3_DATA) && s3_hready)
        m6_s3_req_pend_tmp <= 1'b0;
  end
assign m6_s3_req_pend = m6_s3_req_pend_tmp && (~((m6_cur_st[48:0] == S_S3_DATA) && s3_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m6_s4_req_pend_tmp <= 1'b0;
    else if(m6_latch_cmd && m6_s4_req)
        m6_s4_req_pend_tmp <= 1'b1;
    else if((m6_cur_st[48:0] == S_S4_DATA) && s4_hready)
        m6_s4_req_pend_tmp <= 1'b0;
  end
assign m6_s4_req_pend = m6_s4_req_pend_tmp && (~((m6_cur_st[48:0] == S_S4_DATA) && s4_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m6_s5_req_pend_tmp <= 1'b0;
    else if(m6_latch_cmd && m6_s5_req)
        m6_s5_req_pend_tmp <= 1'b1;
    else if((m6_cur_st[48:0] == S_S5_DATA) && s5_hready)
        m6_s5_req_pend_tmp <= 1'b0;
  end
assign m6_s5_req_pend = m6_s5_req_pend_tmp && (~((m6_cur_st[48:0] == S_S5_DATA) && s5_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m6_s6_req_pend_tmp <= 1'b0;
    else if(m6_latch_cmd && m6_s6_req)
        m6_s6_req_pend_tmp <= 1'b1;
    else if((m6_cur_st[48:0] == S_S6_DATA) && s6_hready)
        m6_s6_req_pend_tmp <= 1'b0;
  end
assign m6_s6_req_pend = m6_s6_req_pend_tmp && (~((m6_cur_st[48:0] == S_S6_DATA) && s6_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m6_s7_req_pend_tmp <= 1'b0;
    else if(m6_latch_cmd && m6_s7_req)
        m6_s7_req_pend_tmp <= 1'b1;
    else if((m6_cur_st[48:0] == S_S7_DATA) && s7_hready)
        m6_s7_req_pend_tmp <= 1'b0;
  end
assign m6_s7_req_pend = m6_s7_req_pend_tmp && (~((m6_cur_st[48:0] == S_S7_DATA) && s7_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m6_s8_req_pend_tmp <= 1'b0;
    else if(m6_latch_cmd && m6_s8_req)
        m6_s8_req_pend_tmp <= 1'b1;
    else if((m6_cur_st[48:0] == S_S8_DATA) && s8_hready)
        m6_s8_req_pend_tmp <= 1'b0;
  end
assign m6_s8_req_pend = m6_s8_req_pend_tmp && (~((m6_cur_st[48:0] == S_S8_DATA) && s8_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m6_s9_req_pend_tmp <= 1'b0;
    else if(m6_latch_cmd && m6_s9_req)
        m6_s9_req_pend_tmp <= 1'b1;
    else if((m6_cur_st[48:0] == S_S9_DATA) && s9_hready)
        m6_s9_req_pend_tmp <= 1'b0;
  end
assign m6_s9_req_pend = m6_s9_req_pend_tmp && (~((m6_cur_st[48:0] == S_S9_DATA) && s9_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m6_s10_req_pend_tmp <= 1'b0;
    else if(m6_latch_cmd && m6_s10_req)
        m6_s10_req_pend_tmp <= 1'b1;
    else if((m6_cur_st[48:0] == S_S10_DATA) && s10_hready)
        m6_s10_req_pend_tmp <= 1'b0;
  end
assign m6_s10_req_pend = m6_s10_req_pend_tmp && (~((m6_cur_st[48:0] == S_S10_DATA) && s10_hready));
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
        m6_s11_req_pend_tmp <= 1'b0;
    else if(m6_latch_cmd && m6_s11_req)
        m6_s11_req_pend_tmp <= 1'b1;
    else if((m6_cur_st[48:0] == S_S11_DATA) && s11_hready)
        m6_s11_req_pend_tmp <= 1'b0;
  end
assign m6_s11_req_pend = m6_s11_req_pend_tmp && (~((m6_cur_st[48:0] == S_S11_DATA) && s11_hready));
assign s0_req_pend[7-1:0] = {
                        m0_s0_req_pend,
                        m1_s0_req_pend,
                        m2_s0_req_pend,
                        m3_s0_req_pend,
                        m4_s0_req_pend,
                        m5_s0_req_pend,
                        m6_s0_req_pend};
assign s1_req_pend[7-1:0] = {
                        m0_s1_req_pend,
                        m1_s1_req_pend,
                        m2_s1_req_pend,
                        m3_s1_req_pend,
                        m4_s1_req_pend,
                        m5_s1_req_pend,
                        m6_s1_req_pend};
assign s2_req_pend[7-1:0] = {
                        m0_s2_req_pend,
                        m1_s2_req_pend,
                        m2_s2_req_pend,
                        m3_s2_req_pend,
                        m4_s2_req_pend,
                        m5_s2_req_pend,
                        m6_s2_req_pend};
assign s3_req_pend[7-1:0] = {
                        m0_s3_req_pend,
                        m1_s3_req_pend,
                        m2_s3_req_pend,
                        m3_s3_req_pend,
                        m4_s3_req_pend,
                        m5_s3_req_pend,
                        m6_s3_req_pend};
assign s4_req_pend[7-1:0] = {
                        m0_s4_req_pend,
                        m1_s4_req_pend,
                        m2_s4_req_pend,
                        m3_s4_req_pend,
                        m4_s4_req_pend,
                        m5_s4_req_pend,
                        m6_s4_req_pend};
assign s5_req_pend[7-1:0] = {
                        m0_s5_req_pend,
                        m1_s5_req_pend,
                        m2_s5_req_pend,
                        m3_s5_req_pend,
                        m4_s5_req_pend,
                        m5_s5_req_pend,
                        m6_s5_req_pend};
assign s6_req_pend[7-1:0] = {
                        m0_s6_req_pend,
                        m1_s6_req_pend,
                        m2_s6_req_pend,
                        m3_s6_req_pend,
                        m4_s6_req_pend,
                        m5_s6_req_pend,
                        m6_s6_req_pend};
assign s7_req_pend[7-1:0] = {
                        m0_s7_req_pend,
                        m1_s7_req_pend,
                        m2_s7_req_pend,
                        m3_s7_req_pend,
                        m4_s7_req_pend,
                        m5_s7_req_pend,
                        m6_s7_req_pend};
assign s8_req_pend[7-1:0] = {
                        m0_s8_req_pend,
                        m1_s8_req_pend,
                        m2_s8_req_pend,
                        m3_s8_req_pend,
                        m4_s8_req_pend,
                        m5_s8_req_pend,
                        m6_s8_req_pend};
assign s9_req_pend[7-1:0] = {
                        m0_s9_req_pend,
                        m1_s9_req_pend,
                        m2_s9_req_pend,
                        m3_s9_req_pend,
                        m4_s9_req_pend,
                        m5_s9_req_pend,
                        m6_s9_req_pend};
assign s10_req_pend[7-1:0] = {
                        m0_s10_req_pend,
                        m1_s10_req_pend,
                        m2_s10_req_pend,
                        m3_s10_req_pend,
                        m4_s10_req_pend,
                        m5_s10_req_pend,
                        m6_s10_req_pend};
assign s11_req_pend[7-1:0] = {
                        m0_s11_req_pend,
                        m1_s11_req_pend,
                        m2_s11_req_pend,
                        m3_s11_req_pend,
                        m4_s11_req_pend,
                        m5_s11_req_pend,
                        m6_s11_req_pend};
always @( s4_hready
       or s10_hready
       or s1_hready
       or s7_hready
       or s5_hready
       or s6_hready
       or s0_hready
       or s8_hready
       or s2_hready
       or s11_hready
       or s3_hready
       or s9_hready
       or m0_cur_st[48:0])
begin
case(m0_cur_st[48:0])
   S_IDLE : m0_nor_hready = 1'b1;
   S_S0_CMD: m0_nor_hready = 1'b0;
   S_S0_GNT: m0_nor_hready = 1'b0;
   S_S0_WAIT : m0_nor_hready = 1'b0;
   S_S1_CMD: m0_nor_hready = 1'b0;
   S_S1_GNT: m0_nor_hready = 1'b0;
   S_S1_WAIT : m0_nor_hready = 1'b0;
   S_S2_CMD: m0_nor_hready = 1'b0;
   S_S2_GNT: m0_nor_hready = 1'b0;
   S_S2_WAIT : m0_nor_hready = 1'b0;
   S_S3_CMD: m0_nor_hready = 1'b0;
   S_S3_GNT: m0_nor_hready = 1'b0;
   S_S3_WAIT : m0_nor_hready = 1'b0;
   S_S4_CMD: m0_nor_hready = 1'b0;
   S_S4_GNT: m0_nor_hready = 1'b0;
   S_S4_WAIT : m0_nor_hready = 1'b0;
   S_S5_CMD: m0_nor_hready = 1'b0;
   S_S5_GNT: m0_nor_hready = 1'b0;
   S_S5_WAIT : m0_nor_hready = 1'b0;
   S_S6_CMD: m0_nor_hready = 1'b0;
   S_S6_GNT: m0_nor_hready = 1'b0;
   S_S6_WAIT : m0_nor_hready = 1'b0;
   S_S7_CMD: m0_nor_hready = 1'b0;
   S_S7_GNT: m0_nor_hready = 1'b0;
   S_S7_WAIT : m0_nor_hready = 1'b0;
   S_S8_CMD: m0_nor_hready = 1'b0;
   S_S8_GNT: m0_nor_hready = 1'b0;
   S_S8_WAIT : m0_nor_hready = 1'b0;
   S_S9_CMD: m0_nor_hready = 1'b0;
   S_S9_GNT: m0_nor_hready = 1'b0;
   S_S9_WAIT : m0_nor_hready = 1'b0;
   S_S10_CMD: m0_nor_hready = 1'b0;
   S_S10_GNT: m0_nor_hready = 1'b0;
   S_S10_WAIT : m0_nor_hready = 1'b0;
   S_S11_CMD: m0_nor_hready = 1'b0;
   S_S11_GNT: m0_nor_hready = 1'b0;
   S_S11_WAIT : m0_nor_hready = 1'b0;
   S_S0_DATA: m0_nor_hready = s0_hready;
   S_S1_DATA: m0_nor_hready = s1_hready;
   S_S2_DATA: m0_nor_hready = s2_hready;
   S_S3_DATA: m0_nor_hready = s3_hready;
   S_S4_DATA: m0_nor_hready = s4_hready;
   S_S5_DATA: m0_nor_hready = s5_hready;
   S_S6_DATA: m0_nor_hready = s6_hready;
   S_S7_DATA: m0_nor_hready = s7_hready;
   S_S8_DATA: m0_nor_hready = s8_hready;
   S_S9_DATA: m0_nor_hready = s9_hready;
   S_S10_DATA: m0_nor_hready = s10_hready;
   S_S11_DATA: m0_nor_hready = s11_hready;
   default: m0_nor_hready = 1'b1;
endcase
end
always @( s4_hready
       or s10_hready
       or s1_hready
       or s7_hready
       or s5_hready
       or s6_hready
       or m1_cur_st[48:0]
       or s0_hready
       or s8_hready
       or s2_hready
       or s11_hready
       or s3_hready
       or s9_hready)
begin
case(m1_cur_st[48:0])
   S_IDLE : m1_nor_hready = 1'b1;
   S_S0_CMD: m1_nor_hready = 1'b0;
   S_S0_GNT: m1_nor_hready = 1'b0;
   S_S0_WAIT : m1_nor_hready = 1'b0;
   S_S1_CMD: m1_nor_hready = 1'b0;
   S_S1_GNT: m1_nor_hready = 1'b0;
   S_S1_WAIT : m1_nor_hready = 1'b0;
   S_S2_CMD: m1_nor_hready = 1'b0;
   S_S2_GNT: m1_nor_hready = 1'b0;
   S_S2_WAIT : m1_nor_hready = 1'b0;
   S_S3_CMD: m1_nor_hready = 1'b0;
   S_S3_GNT: m1_nor_hready = 1'b0;
   S_S3_WAIT : m1_nor_hready = 1'b0;
   S_S4_CMD: m1_nor_hready = 1'b0;
   S_S4_GNT: m1_nor_hready = 1'b0;
   S_S4_WAIT : m1_nor_hready = 1'b0;
   S_S5_CMD: m1_nor_hready = 1'b0;
   S_S5_GNT: m1_nor_hready = 1'b0;
   S_S5_WAIT : m1_nor_hready = 1'b0;
   S_S6_CMD: m1_nor_hready = 1'b0;
   S_S6_GNT: m1_nor_hready = 1'b0;
   S_S6_WAIT : m1_nor_hready = 1'b0;
   S_S7_CMD: m1_nor_hready = 1'b0;
   S_S7_GNT: m1_nor_hready = 1'b0;
   S_S7_WAIT : m1_nor_hready = 1'b0;
   S_S8_CMD: m1_nor_hready = 1'b0;
   S_S8_GNT: m1_nor_hready = 1'b0;
   S_S8_WAIT : m1_nor_hready = 1'b0;
   S_S9_CMD: m1_nor_hready = 1'b0;
   S_S9_GNT: m1_nor_hready = 1'b0;
   S_S9_WAIT : m1_nor_hready = 1'b0;
   S_S10_CMD: m1_nor_hready = 1'b0;
   S_S10_GNT: m1_nor_hready = 1'b0;
   S_S10_WAIT : m1_nor_hready = 1'b0;
   S_S11_CMD: m1_nor_hready = 1'b0;
   S_S11_GNT: m1_nor_hready = 1'b0;
   S_S11_WAIT : m1_nor_hready = 1'b0;
   S_S0_DATA: m1_nor_hready = s0_hready;
   S_S1_DATA: m1_nor_hready = s1_hready;
   S_S2_DATA: m1_nor_hready = s2_hready;
   S_S3_DATA: m1_nor_hready = s3_hready;
   S_S4_DATA: m1_nor_hready = s4_hready;
   S_S5_DATA: m1_nor_hready = s5_hready;
   S_S6_DATA: m1_nor_hready = s6_hready;
   S_S7_DATA: m1_nor_hready = s7_hready;
   S_S8_DATA: m1_nor_hready = s8_hready;
   S_S9_DATA: m1_nor_hready = s9_hready;
   S_S10_DATA: m1_nor_hready = s10_hready;
   S_S11_DATA: m1_nor_hready = s11_hready;
   default: m1_nor_hready = 1'b1;
endcase
end
always @( s4_hready
       or s10_hready
       or s1_hready
       or s7_hready
       or m2_cur_st[48:0]
       or s5_hready
       or s6_hready
       or s0_hready
       or s8_hready
       or s2_hready
       or s11_hready
       or s3_hready
       or s9_hready)
begin
case(m2_cur_st[48:0])
   S_IDLE : m2_nor_hready = 1'b1;
   S_S0_CMD: m2_nor_hready = 1'b0;
   S_S0_GNT: m2_nor_hready = 1'b0;
   S_S0_WAIT : m2_nor_hready = 1'b0;
   S_S1_CMD: m2_nor_hready = 1'b0;
   S_S1_GNT: m2_nor_hready = 1'b0;
   S_S1_WAIT : m2_nor_hready = 1'b0;
   S_S2_CMD: m2_nor_hready = 1'b0;
   S_S2_GNT: m2_nor_hready = 1'b0;
   S_S2_WAIT : m2_nor_hready = 1'b0;
   S_S3_CMD: m2_nor_hready = 1'b0;
   S_S3_GNT: m2_nor_hready = 1'b0;
   S_S3_WAIT : m2_nor_hready = 1'b0;
   S_S4_CMD: m2_nor_hready = 1'b0;
   S_S4_GNT: m2_nor_hready = 1'b0;
   S_S4_WAIT : m2_nor_hready = 1'b0;
   S_S5_CMD: m2_nor_hready = 1'b0;
   S_S5_GNT: m2_nor_hready = 1'b0;
   S_S5_WAIT : m2_nor_hready = 1'b0;
   S_S6_CMD: m2_nor_hready = 1'b0;
   S_S6_GNT: m2_nor_hready = 1'b0;
   S_S6_WAIT : m2_nor_hready = 1'b0;
   S_S7_CMD: m2_nor_hready = 1'b0;
   S_S7_GNT: m2_nor_hready = 1'b0;
   S_S7_WAIT : m2_nor_hready = 1'b0;
   S_S8_CMD: m2_nor_hready = 1'b0;
   S_S8_GNT: m2_nor_hready = 1'b0;
   S_S8_WAIT : m2_nor_hready = 1'b0;
   S_S9_CMD: m2_nor_hready = 1'b0;
   S_S9_GNT: m2_nor_hready = 1'b0;
   S_S9_WAIT : m2_nor_hready = 1'b0;
   S_S10_CMD: m2_nor_hready = 1'b0;
   S_S10_GNT: m2_nor_hready = 1'b0;
   S_S10_WAIT : m2_nor_hready = 1'b0;
   S_S11_CMD: m2_nor_hready = 1'b0;
   S_S11_GNT: m2_nor_hready = 1'b0;
   S_S11_WAIT : m2_nor_hready = 1'b0;
   S_S0_DATA: m2_nor_hready = s0_hready;
   S_S1_DATA: m2_nor_hready = s1_hready;
   S_S2_DATA: m2_nor_hready = s2_hready;
   S_S3_DATA: m2_nor_hready = s3_hready;
   S_S4_DATA: m2_nor_hready = s4_hready;
   S_S5_DATA: m2_nor_hready = s5_hready;
   S_S6_DATA: m2_nor_hready = s6_hready;
   S_S7_DATA: m2_nor_hready = s7_hready;
   S_S8_DATA: m2_nor_hready = s8_hready;
   S_S9_DATA: m2_nor_hready = s9_hready;
   S_S10_DATA: m2_nor_hready = s10_hready;
   S_S11_DATA: m2_nor_hready = s11_hready;
   default: m2_nor_hready = 1'b1;
endcase
end
always @( s4_hready
       or s10_hready
       or s1_hready
       or s7_hready
       or s5_hready
       or s6_hready
       or s0_hready
       or s8_hready
       or m3_cur_st[48:0]
       or s2_hready
       or s11_hready
       or s3_hready
       or s9_hready)
begin
case(m3_cur_st[48:0])
   S_IDLE : m3_nor_hready = 1'b1;
   S_S0_CMD: m3_nor_hready = 1'b0;
   S_S0_GNT: m3_nor_hready = 1'b0;
   S_S0_WAIT : m3_nor_hready = 1'b0;
   S_S1_CMD: m3_nor_hready = 1'b0;
   S_S1_GNT: m3_nor_hready = 1'b0;
   S_S1_WAIT : m3_nor_hready = 1'b0;
   S_S2_CMD: m3_nor_hready = 1'b0;
   S_S2_GNT: m3_nor_hready = 1'b0;
   S_S2_WAIT : m3_nor_hready = 1'b0;
   S_S3_CMD: m3_nor_hready = 1'b0;
   S_S3_GNT: m3_nor_hready = 1'b0;
   S_S3_WAIT : m3_nor_hready = 1'b0;
   S_S4_CMD: m3_nor_hready = 1'b0;
   S_S4_GNT: m3_nor_hready = 1'b0;
   S_S4_WAIT : m3_nor_hready = 1'b0;
   S_S5_CMD: m3_nor_hready = 1'b0;
   S_S5_GNT: m3_nor_hready = 1'b0;
   S_S5_WAIT : m3_nor_hready = 1'b0;
   S_S6_CMD: m3_nor_hready = 1'b0;
   S_S6_GNT: m3_nor_hready = 1'b0;
   S_S6_WAIT : m3_nor_hready = 1'b0;
   S_S7_CMD: m3_nor_hready = 1'b0;
   S_S7_GNT: m3_nor_hready = 1'b0;
   S_S7_WAIT : m3_nor_hready = 1'b0;
   S_S8_CMD: m3_nor_hready = 1'b0;
   S_S8_GNT: m3_nor_hready = 1'b0;
   S_S8_WAIT : m3_nor_hready = 1'b0;
   S_S9_CMD: m3_nor_hready = 1'b0;
   S_S9_GNT: m3_nor_hready = 1'b0;
   S_S9_WAIT : m3_nor_hready = 1'b0;
   S_S10_CMD: m3_nor_hready = 1'b0;
   S_S10_GNT: m3_nor_hready = 1'b0;
   S_S10_WAIT : m3_nor_hready = 1'b0;
   S_S11_CMD: m3_nor_hready = 1'b0;
   S_S11_GNT: m3_nor_hready = 1'b0;
   S_S11_WAIT : m3_nor_hready = 1'b0;
   S_S0_DATA: m3_nor_hready = s0_hready;
   S_S1_DATA: m3_nor_hready = s1_hready;
   S_S2_DATA: m3_nor_hready = s2_hready;
   S_S3_DATA: m3_nor_hready = s3_hready;
   S_S4_DATA: m3_nor_hready = s4_hready;
   S_S5_DATA: m3_nor_hready = s5_hready;
   S_S6_DATA: m3_nor_hready = s6_hready;
   S_S7_DATA: m3_nor_hready = s7_hready;
   S_S8_DATA: m3_nor_hready = s8_hready;
   S_S9_DATA: m3_nor_hready = s9_hready;
   S_S10_DATA: m3_nor_hready = s10_hready;
   S_S11_DATA: m3_nor_hready = s11_hready;
   default: m3_nor_hready = 1'b1;
endcase
end
always @( s4_hready
       or s10_hready
       or s1_hready
       or s7_hready
       or s5_hready
       or s6_hready
       or s0_hready
       or s8_hready
       or s2_hready
       or s11_hready
       or m4_cur_st[48:0]
       or s3_hready
       or s9_hready)
begin
case(m4_cur_st[48:0])
   S_IDLE : m4_nor_hready = 1'b1;
   S_S0_CMD: m4_nor_hready = 1'b0;
   S_S0_GNT: m4_nor_hready = 1'b0;
   S_S0_WAIT : m4_nor_hready = 1'b0;
   S_S1_CMD: m4_nor_hready = 1'b0;
   S_S1_GNT: m4_nor_hready = 1'b0;
   S_S1_WAIT : m4_nor_hready = 1'b0;
   S_S2_CMD: m4_nor_hready = 1'b0;
   S_S2_GNT: m4_nor_hready = 1'b0;
   S_S2_WAIT : m4_nor_hready = 1'b0;
   S_S3_CMD: m4_nor_hready = 1'b0;
   S_S3_GNT: m4_nor_hready = 1'b0;
   S_S3_WAIT : m4_nor_hready = 1'b0;
   S_S4_CMD: m4_nor_hready = 1'b0;
   S_S4_GNT: m4_nor_hready = 1'b0;
   S_S4_WAIT : m4_nor_hready = 1'b0;
   S_S5_CMD: m4_nor_hready = 1'b0;
   S_S5_GNT: m4_nor_hready = 1'b0;
   S_S5_WAIT : m4_nor_hready = 1'b0;
   S_S6_CMD: m4_nor_hready = 1'b0;
   S_S6_GNT: m4_nor_hready = 1'b0;
   S_S6_WAIT : m4_nor_hready = 1'b0;
   S_S7_CMD: m4_nor_hready = 1'b0;
   S_S7_GNT: m4_nor_hready = 1'b0;
   S_S7_WAIT : m4_nor_hready = 1'b0;
   S_S8_CMD: m4_nor_hready = 1'b0;
   S_S8_GNT: m4_nor_hready = 1'b0;
   S_S8_WAIT : m4_nor_hready = 1'b0;
   S_S9_CMD: m4_nor_hready = 1'b0;
   S_S9_GNT: m4_nor_hready = 1'b0;
   S_S9_WAIT : m4_nor_hready = 1'b0;
   S_S10_CMD: m4_nor_hready = 1'b0;
   S_S10_GNT: m4_nor_hready = 1'b0;
   S_S10_WAIT : m4_nor_hready = 1'b0;
   S_S11_CMD: m4_nor_hready = 1'b0;
   S_S11_GNT: m4_nor_hready = 1'b0;
   S_S11_WAIT : m4_nor_hready = 1'b0;
   S_S0_DATA: m4_nor_hready = s0_hready;
   S_S1_DATA: m4_nor_hready = s1_hready;
   S_S2_DATA: m4_nor_hready = s2_hready;
   S_S3_DATA: m4_nor_hready = s3_hready;
   S_S4_DATA: m4_nor_hready = s4_hready;
   S_S5_DATA: m4_nor_hready = s5_hready;
   S_S6_DATA: m4_nor_hready = s6_hready;
   S_S7_DATA: m4_nor_hready = s7_hready;
   S_S8_DATA: m4_nor_hready = s8_hready;
   S_S9_DATA: m4_nor_hready = s9_hready;
   S_S10_DATA: m4_nor_hready = s10_hready;
   S_S11_DATA: m4_nor_hready = s11_hready;
   default: m4_nor_hready = 1'b1;
endcase
end
always @( s4_hready
       or s10_hready
       or s1_hready
       or s7_hready
       or s5_hready
       or s6_hready
       or s0_hready
       or s8_hready
       or m5_cur_st[48:0]
       or s2_hready
       or s11_hready
       or s3_hready
       or s9_hready)
begin
case(m5_cur_st[48:0])
   S_IDLE : m5_nor_hready = 1'b1;
   S_S0_CMD: m5_nor_hready = 1'b0;
   S_S0_GNT: m5_nor_hready = 1'b0;
   S_S0_WAIT : m5_nor_hready = 1'b0;
   S_S1_CMD: m5_nor_hready = 1'b0;
   S_S1_GNT: m5_nor_hready = 1'b0;
   S_S1_WAIT : m5_nor_hready = 1'b0;
   S_S2_CMD: m5_nor_hready = 1'b0;
   S_S2_GNT: m5_nor_hready = 1'b0;
   S_S2_WAIT : m5_nor_hready = 1'b0;
   S_S3_CMD: m5_nor_hready = 1'b0;
   S_S3_GNT: m5_nor_hready = 1'b0;
   S_S3_WAIT : m5_nor_hready = 1'b0;
   S_S4_CMD: m5_nor_hready = 1'b0;
   S_S4_GNT: m5_nor_hready = 1'b0;
   S_S4_WAIT : m5_nor_hready = 1'b0;
   S_S5_CMD: m5_nor_hready = 1'b0;
   S_S5_GNT: m5_nor_hready = 1'b0;
   S_S5_WAIT : m5_nor_hready = 1'b0;
   S_S6_CMD: m5_nor_hready = 1'b0;
   S_S6_GNT: m5_nor_hready = 1'b0;
   S_S6_WAIT : m5_nor_hready = 1'b0;
   S_S7_CMD: m5_nor_hready = 1'b0;
   S_S7_GNT: m5_nor_hready = 1'b0;
   S_S7_WAIT : m5_nor_hready = 1'b0;
   S_S8_CMD: m5_nor_hready = 1'b0;
   S_S8_GNT: m5_nor_hready = 1'b0;
   S_S8_WAIT : m5_nor_hready = 1'b0;
   S_S9_CMD: m5_nor_hready = 1'b0;
   S_S9_GNT: m5_nor_hready = 1'b0;
   S_S9_WAIT : m5_nor_hready = 1'b0;
   S_S10_CMD: m5_nor_hready = 1'b0;
   S_S10_GNT: m5_nor_hready = 1'b0;
   S_S10_WAIT : m5_nor_hready = 1'b0;
   S_S11_CMD: m5_nor_hready = 1'b0;
   S_S11_GNT: m5_nor_hready = 1'b0;
   S_S11_WAIT : m5_nor_hready = 1'b0;
   S_S0_DATA: m5_nor_hready = s0_hready;
   S_S1_DATA: m5_nor_hready = s1_hready;
   S_S2_DATA: m5_nor_hready = s2_hready;
   S_S3_DATA: m5_nor_hready = s3_hready;
   S_S4_DATA: m5_nor_hready = s4_hready;
   S_S5_DATA: m5_nor_hready = s5_hready;
   S_S6_DATA: m5_nor_hready = s6_hready;
   S_S7_DATA: m5_nor_hready = s7_hready;
   S_S8_DATA: m5_nor_hready = s8_hready;
   S_S9_DATA: m5_nor_hready = s9_hready;
   S_S10_DATA: m5_nor_hready = s10_hready;
   S_S11_DATA: m5_nor_hready = s11_hready;
   default: m5_nor_hready = 1'b1;
endcase
end
always @( s4_hready
       or s10_hready
       or s1_hready
       or s7_hready
       or s5_hready
       or s6_hready
       or m6_cur_st[48:0]
       or s0_hready
       or s8_hready
       or s2_hready
       or s11_hready
       or s3_hready
       or s9_hready)
begin
case(m6_cur_st[48:0])
   S_IDLE : m6_nor_hready = 1'b1;
   S_S0_CMD: m6_nor_hready = 1'b0;
   S_S0_GNT: m6_nor_hready = 1'b0;
   S_S0_WAIT : m6_nor_hready = 1'b0;
   S_S1_CMD: m6_nor_hready = 1'b0;
   S_S1_GNT: m6_nor_hready = 1'b0;
   S_S1_WAIT : m6_nor_hready = 1'b0;
   S_S2_CMD: m6_nor_hready = 1'b0;
   S_S2_GNT: m6_nor_hready = 1'b0;
   S_S2_WAIT : m6_nor_hready = 1'b0;
   S_S3_CMD: m6_nor_hready = 1'b0;
   S_S3_GNT: m6_nor_hready = 1'b0;
   S_S3_WAIT : m6_nor_hready = 1'b0;
   S_S4_CMD: m6_nor_hready = 1'b0;
   S_S4_GNT: m6_nor_hready = 1'b0;
   S_S4_WAIT : m6_nor_hready = 1'b0;
   S_S5_CMD: m6_nor_hready = 1'b0;
   S_S5_GNT: m6_nor_hready = 1'b0;
   S_S5_WAIT : m6_nor_hready = 1'b0;
   S_S6_CMD: m6_nor_hready = 1'b0;
   S_S6_GNT: m6_nor_hready = 1'b0;
   S_S6_WAIT : m6_nor_hready = 1'b0;
   S_S7_CMD: m6_nor_hready = 1'b0;
   S_S7_GNT: m6_nor_hready = 1'b0;
   S_S7_WAIT : m6_nor_hready = 1'b0;
   S_S8_CMD: m6_nor_hready = 1'b0;
   S_S8_GNT: m6_nor_hready = 1'b0;
   S_S8_WAIT : m6_nor_hready = 1'b0;
   S_S9_CMD: m6_nor_hready = 1'b0;
   S_S9_GNT: m6_nor_hready = 1'b0;
   S_S9_WAIT : m6_nor_hready = 1'b0;
   S_S10_CMD: m6_nor_hready = 1'b0;
   S_S10_GNT: m6_nor_hready = 1'b0;
   S_S10_WAIT : m6_nor_hready = 1'b0;
   S_S11_CMD: m6_nor_hready = 1'b0;
   S_S11_GNT: m6_nor_hready = 1'b0;
   S_S11_WAIT : m6_nor_hready = 1'b0;
   S_S0_DATA: m6_nor_hready = s0_hready;
   S_S1_DATA: m6_nor_hready = s1_hready;
   S_S2_DATA: m6_nor_hready = s2_hready;
   S_S3_DATA: m6_nor_hready = s3_hready;
   S_S4_DATA: m6_nor_hready = s4_hready;
   S_S5_DATA: m6_nor_hready = s5_hready;
   S_S6_DATA: m6_nor_hready = s6_hready;
   S_S7_DATA: m6_nor_hready = s7_hready;
   S_S8_DATA: m6_nor_hready = s8_hready;
   S_S9_DATA: m6_nor_hready = s9_hready;
   S_S10_DATA: m6_nor_hready = s10_hready;
   S_S11_DATA: m6_nor_hready = s11_hready;
   default: m6_nor_hready = 1'b1;
endcase
end
endmodule
module ahb_matrix_7_12_dec(
  hclk,
  hresetn,
  m0_haddr,
  m0_hburst,
  m0_hgrant,
  m0_hprot,
  m0_hrdata,
  m0_hready,
  m0_hresp,
  m0_hsize,
  m0_htrans,
  m0_hwdata,
  m0_hwrite,
  m0_latch_cmd,
  m0_nor_hready,
  m0_s0_cmd_cur,
  m0_s0_cmd_last,
  m0_s0_data,
  m0_s0_req,
  m0_s10_cmd_cur,
  m0_s10_cmd_last,
  m0_s10_data,
  m0_s10_req,
  m0_s11_cmd_cur,
  m0_s11_cmd_last,
  m0_s11_data,
  m0_s11_req,
  m0_s1_cmd_cur,
  m0_s1_cmd_last,
  m0_s1_data,
  m0_s1_req,
  m0_s2_cmd_cur,
  m0_s2_cmd_last,
  m0_s2_data,
  m0_s2_req,
  m0_s3_cmd_cur,
  m0_s3_cmd_last,
  m0_s3_data,
  m0_s3_req,
  m0_s4_cmd_cur,
  m0_s4_cmd_last,
  m0_s4_data,
  m0_s4_req,
  m0_s5_cmd_cur,
  m0_s5_cmd_last,
  m0_s5_data,
  m0_s5_req,
  m0_s6_cmd_cur,
  m0_s6_cmd_last,
  m0_s6_data,
  m0_s6_req,
  m0_s7_cmd_cur,
  m0_s7_cmd_last,
  m0_s7_data,
  m0_s7_req,
  m0_s8_cmd_cur,
  m0_s8_cmd_last,
  m0_s8_data,
  m0_s8_req,
  m0_s9_cmd_cur,
  m0_s9_cmd_last,
  m0_s9_data,
  m0_s9_req,
  m1_haddr,
  m1_hburst,
  m1_hgrant,
  m1_hprot,
  m1_hrdata,
  m1_hready,
  m1_hresp,
  m1_hsize,
  m1_htrans,
  m1_hwdata,
  m1_hwrite,
  m1_latch_cmd,
  m1_nor_hready,
  m1_s0_cmd_cur,
  m1_s0_cmd_last,
  m1_s0_data,
  m1_s0_req,
  m1_s10_cmd_cur,
  m1_s10_cmd_last,
  m1_s10_data,
  m1_s10_req,
  m1_s11_cmd_cur,
  m1_s11_cmd_last,
  m1_s11_data,
  m1_s11_req,
  m1_s1_cmd_cur,
  m1_s1_cmd_last,
  m1_s1_data,
  m1_s1_req,
  m1_s2_cmd_cur,
  m1_s2_cmd_last,
  m1_s2_data,
  m1_s2_req,
  m1_s3_cmd_cur,
  m1_s3_cmd_last,
  m1_s3_data,
  m1_s3_req,
  m1_s4_cmd_cur,
  m1_s4_cmd_last,
  m1_s4_data,
  m1_s4_req,
  m1_s5_cmd_cur,
  m1_s5_cmd_last,
  m1_s5_data,
  m1_s5_req,
  m1_s6_cmd_cur,
  m1_s6_cmd_last,
  m1_s6_data,
  m1_s6_req,
  m1_s7_cmd_cur,
  m1_s7_cmd_last,
  m1_s7_data,
  m1_s7_req,
  m1_s8_cmd_cur,
  m1_s8_cmd_last,
  m1_s8_data,
  m1_s8_req,
  m1_s9_cmd_cur,
  m1_s9_cmd_last,
  m1_s9_data,
  m1_s9_req,
  m2_haddr,
  m2_hburst,
  m2_hgrant,
  m2_hprot,
  m2_hrdata,
  m2_hready,
  m2_hresp,
  m2_hsize,
  m2_htrans,
  m2_hwdata,
  m2_hwrite,
  m2_latch_cmd,
  m2_nor_hready,
  m2_s0_cmd_cur,
  m2_s0_cmd_last,
  m2_s0_data,
  m2_s0_req,
  m2_s10_cmd_cur,
  m2_s10_cmd_last,
  m2_s10_data,
  m2_s10_req,
  m2_s11_cmd_cur,
  m2_s11_cmd_last,
  m2_s11_data,
  m2_s11_req,
  m2_s1_cmd_cur,
  m2_s1_cmd_last,
  m2_s1_data,
  m2_s1_req,
  m2_s2_cmd_cur,
  m2_s2_cmd_last,
  m2_s2_data,
  m2_s2_req,
  m2_s3_cmd_cur,
  m2_s3_cmd_last,
  m2_s3_data,
  m2_s3_req,
  m2_s4_cmd_cur,
  m2_s4_cmd_last,
  m2_s4_data,
  m2_s4_req,
  m2_s5_cmd_cur,
  m2_s5_cmd_last,
  m2_s5_data,
  m2_s5_req,
  m2_s6_cmd_cur,
  m2_s6_cmd_last,
  m2_s6_data,
  m2_s6_req,
  m2_s7_cmd_cur,
  m2_s7_cmd_last,
  m2_s7_data,
  m2_s7_req,
  m2_s8_cmd_cur,
  m2_s8_cmd_last,
  m2_s8_data,
  m2_s8_req,
  m2_s9_cmd_cur,
  m2_s9_cmd_last,
  m2_s9_data,
  m2_s9_req,
  m3_haddr,
  m3_hburst,
  m3_hgrant,
  m3_hprot,
  m3_hrdata,
  m3_hready,
  m3_hresp,
  m3_hsize,
  m3_htrans,
  m3_hwdata,
  m3_hwrite,
  m3_latch_cmd,
  m3_nor_hready,
  m3_s0_cmd_cur,
  m3_s0_cmd_last,
  m3_s0_data,
  m3_s0_req,
  m3_s10_cmd_cur,
  m3_s10_cmd_last,
  m3_s10_data,
  m3_s10_req,
  m3_s11_cmd_cur,
  m3_s11_cmd_last,
  m3_s11_data,
  m3_s11_req,
  m3_s1_cmd_cur,
  m3_s1_cmd_last,
  m3_s1_data,
  m3_s1_req,
  m3_s2_cmd_cur,
  m3_s2_cmd_last,
  m3_s2_data,
  m3_s2_req,
  m3_s3_cmd_cur,
  m3_s3_cmd_last,
  m3_s3_data,
  m3_s3_req,
  m3_s4_cmd_cur,
  m3_s4_cmd_last,
  m3_s4_data,
  m3_s4_req,
  m3_s5_cmd_cur,
  m3_s5_cmd_last,
  m3_s5_data,
  m3_s5_req,
  m3_s6_cmd_cur,
  m3_s6_cmd_last,
  m3_s6_data,
  m3_s6_req,
  m3_s7_cmd_cur,
  m3_s7_cmd_last,
  m3_s7_data,
  m3_s7_req,
  m3_s8_cmd_cur,
  m3_s8_cmd_last,
  m3_s8_data,
  m3_s8_req,
  m3_s9_cmd_cur,
  m3_s9_cmd_last,
  m3_s9_data,
  m3_s9_req,
  m4_haddr,
  m4_hburst,
  m4_hgrant,
  m4_hprot,
  m4_hrdata,
  m4_hready,
  m4_hresp,
  m4_hsize,
  m4_htrans,
  m4_hwdata,
  m4_hwrite,
  m4_latch_cmd,
  m4_nor_hready,
  m4_s0_cmd_cur,
  m4_s0_cmd_last,
  m4_s0_data,
  m4_s0_req,
  m4_s10_cmd_cur,
  m4_s10_cmd_last,
  m4_s10_data,
  m4_s10_req,
  m4_s11_cmd_cur,
  m4_s11_cmd_last,
  m4_s11_data,
  m4_s11_req,
  m4_s1_cmd_cur,
  m4_s1_cmd_last,
  m4_s1_data,
  m4_s1_req,
  m4_s2_cmd_cur,
  m4_s2_cmd_last,
  m4_s2_data,
  m4_s2_req,
  m4_s3_cmd_cur,
  m4_s3_cmd_last,
  m4_s3_data,
  m4_s3_req,
  m4_s4_cmd_cur,
  m4_s4_cmd_last,
  m4_s4_data,
  m4_s4_req,
  m4_s5_cmd_cur,
  m4_s5_cmd_last,
  m4_s5_data,
  m4_s5_req,
  m4_s6_cmd_cur,
  m4_s6_cmd_last,
  m4_s6_data,
  m4_s6_req,
  m4_s7_cmd_cur,
  m4_s7_cmd_last,
  m4_s7_data,
  m4_s7_req,
  m4_s8_cmd_cur,
  m4_s8_cmd_last,
  m4_s8_data,
  m4_s8_req,
  m4_s9_cmd_cur,
  m4_s9_cmd_last,
  m4_s9_data,
  m4_s9_req,
  m5_haddr,
  m5_hburst,
  m5_hgrant,
  m5_hprot,
  m5_hrdata,
  m5_hready,
  m5_hresp,
  m5_hsize,
  m5_htrans,
  m5_hwdata,
  m5_hwrite,
  m5_latch_cmd,
  m5_nor_hready,
  m5_s0_cmd_cur,
  m5_s0_cmd_last,
  m5_s0_data,
  m5_s0_req,
  m5_s10_cmd_cur,
  m5_s10_cmd_last,
  m5_s10_data,
  m5_s10_req,
  m5_s11_cmd_cur,
  m5_s11_cmd_last,
  m5_s11_data,
  m5_s11_req,
  m5_s1_cmd_cur,
  m5_s1_cmd_last,
  m5_s1_data,
  m5_s1_req,
  m5_s2_cmd_cur,
  m5_s2_cmd_last,
  m5_s2_data,
  m5_s2_req,
  m5_s3_cmd_cur,
  m5_s3_cmd_last,
  m5_s3_data,
  m5_s3_req,
  m5_s4_cmd_cur,
  m5_s4_cmd_last,
  m5_s4_data,
  m5_s4_req,
  m5_s5_cmd_cur,
  m5_s5_cmd_last,
  m5_s5_data,
  m5_s5_req,
  m5_s6_cmd_cur,
  m5_s6_cmd_last,
  m5_s6_data,
  m5_s6_req,
  m5_s7_cmd_cur,
  m5_s7_cmd_last,
  m5_s7_data,
  m5_s7_req,
  m5_s8_cmd_cur,
  m5_s8_cmd_last,
  m5_s8_data,
  m5_s8_req,
  m5_s9_cmd_cur,
  m5_s9_cmd_last,
  m5_s9_data,
  m5_s9_req,
  m6_haddr,
  m6_hburst,
  m6_hgrant,
  m6_hprot,
  m6_hrdata,
  m6_hready,
  m6_hresp,
  m6_hsize,
  m6_htrans,
  m6_hwdata,
  m6_hwrite,
  m6_latch_cmd,
  m6_nor_hready,
  m6_s0_cmd_cur,
  m6_s0_cmd_last,
  m6_s0_data,
  m6_s0_req,
  m6_s10_cmd_cur,
  m6_s10_cmd_last,
  m6_s10_data,
  m6_s10_req,
  m6_s11_cmd_cur,
  m6_s11_cmd_last,
  m6_s11_data,
  m6_s11_req,
  m6_s1_cmd_cur,
  m6_s1_cmd_last,
  m6_s1_data,
  m6_s1_req,
  m6_s2_cmd_cur,
  m6_s2_cmd_last,
  m6_s2_data,
  m6_s2_req,
  m6_s3_cmd_cur,
  m6_s3_cmd_last,
  m6_s3_data,
  m6_s3_req,
  m6_s4_cmd_cur,
  m6_s4_cmd_last,
  m6_s4_data,
  m6_s4_req,
  m6_s5_cmd_cur,
  m6_s5_cmd_last,
  m6_s5_data,
  m6_s5_req,
  m6_s6_cmd_cur,
  m6_s6_cmd_last,
  m6_s6_data,
  m6_s6_req,
  m6_s7_cmd_cur,
  m6_s7_cmd_last,
  m6_s7_data,
  m6_s7_req,
  m6_s8_cmd_cur,
  m6_s8_cmd_last,
  m6_s8_data,
  m6_s8_req,
  m6_s9_cmd_cur,
  m6_s9_cmd_last,
  m6_s9_data,
  m6_s9_req,
  s0_haddr,
  s0_hburst,
  s0_hprot,
  s0_hrdata,
  s0_hresp,
  s0_hselx,
  s0_hsize,
  s0_htrans,
  s0_hwdata,
  s0_hwrite,
  s0_req,
  s10_haddr,
  s10_hburst,
  s10_hprot,
  s10_hrdata,
  s10_hresp,
  s10_hselx,
  s10_hsize,
  s10_htrans,
  s10_hwdata,
  s10_hwrite,
  s10_req,
  s11_haddr,
  s11_hburst,
  s11_hprot,
  s11_hrdata,
  s11_hresp,
  s11_hselx,
  s11_hsize,
  s11_htrans,
  s11_hwdata,
  s11_hwrite,
  s11_req,
  s1_haddr,
  s1_hburst,
  s1_hprot,
  s1_hrdata,
  s1_hresp,
  s1_hselx,
  s1_hsize,
  s1_htrans,
  s1_hwdata,
  s1_hwrite,
  s1_req,
  s2_haddr,
  s2_hburst,
  s2_hprot,
  s2_hrdata,
  s2_hresp,
  s2_hselx,
  s2_hsize,
  s2_htrans,
  s2_hwdata,
  s2_hwrite,
  s2_req,
  s3_haddr,
  s3_hburst,
  s3_hprot,
  s3_hrdata,
  s3_hresp,
  s3_hselx,
  s3_hsize,
  s3_htrans,
  s3_hwdata,
  s3_hwrite,
  s3_req,
  s4_haddr,
  s4_hburst,
  s4_hprot,
  s4_hrdata,
  s4_hresp,
  s4_hselx,
  s4_hsize,
  s4_htrans,
  s4_hwdata,
  s4_hwrite,
  s4_req,
  s5_haddr,
  s5_hburst,
  s5_hprot,
  s5_hrdata,
  s5_hresp,
  s5_hselx,
  s5_hsize,
  s5_htrans,
  s5_hwdata,
  s5_hwrite,
  s5_req,
  s6_haddr,
  s6_hburst,
  s6_hprot,
  s6_hrdata,
  s6_hresp,
  s6_hselx,
  s6_hsize,
  s6_htrans,
  s6_hwdata,
  s6_hwrite,
  s6_req,
  s7_haddr,
  s7_hburst,
  s7_hprot,
  s7_hrdata,
  s7_hresp,
  s7_hselx,
  s7_hsize,
  s7_htrans,
  s7_hwdata,
  s7_hwrite,
  s7_req,
  s8_haddr,
  s8_hburst,
  s8_hprot,
  s8_hrdata,
  s8_hresp,
  s8_hselx,
  s8_hsize,
  s8_htrans,
  s8_hwdata,
  s8_hwrite,
  s8_req,
  s9_haddr,
  s9_hburst,
  s9_hprot,
  s9_hrdata,
  s9_hresp,
  s9_hselx,
  s9_hsize,
  s9_htrans,
  s9_hwdata,
  s9_hwrite,
  s9_req
);
input           hclk;           
input           hresetn;        
input   [31:0]  m0_haddr;       
input   [2 :0]  m0_hburst;      
input   [3 :0]  m0_hprot;       
input   [2 :0]  m0_hsize;       
input   [1 :0]  m0_htrans;      
input   [31:0]  m0_hwdata;      
input           m0_hwrite;      
input           m0_latch_cmd;   
input           m0_nor_hready;  
input           m0_s0_cmd_cur;  
input           m0_s0_cmd_last; 
input           m0_s0_data;     
input           m0_s10_cmd_cur; 
input           m0_s10_cmd_last; 
input           m0_s10_data;    
input           m0_s11_cmd_cur; 
input           m0_s11_cmd_last; 
input           m0_s11_data;    
input           m0_s1_cmd_cur;  
input           m0_s1_cmd_last; 
input           m0_s1_data;     
input           m0_s2_cmd_cur;  
input           m0_s2_cmd_last; 
input           m0_s2_data;     
input           m0_s3_cmd_cur;  
input           m0_s3_cmd_last; 
input           m0_s3_data;     
input           m0_s4_cmd_cur;  
input           m0_s4_cmd_last; 
input           m0_s4_data;     
input           m0_s5_cmd_cur;  
input           m0_s5_cmd_last; 
input           m0_s5_data;     
input           m0_s6_cmd_cur;  
input           m0_s6_cmd_last; 
input           m0_s6_data;     
input           m0_s7_cmd_cur;  
input           m0_s7_cmd_last; 
input           m0_s7_data;     
input           m0_s8_cmd_cur;  
input           m0_s8_cmd_last; 
input           m0_s8_data;     
input           m0_s9_cmd_cur;  
input           m0_s9_cmd_last; 
input           m0_s9_data;     
input   [31:0]  m1_haddr;       
input   [2 :0]  m1_hburst;      
input   [3 :0]  m1_hprot;       
input   [2 :0]  m1_hsize;       
input   [1 :0]  m1_htrans;      
input   [31:0]  m1_hwdata;      
input           m1_hwrite;      
input           m1_latch_cmd;   
input           m1_nor_hready;  
input           m1_s0_cmd_cur;  
input           m1_s0_cmd_last; 
input           m1_s0_data;     
input           m1_s10_cmd_cur; 
input           m1_s10_cmd_last; 
input           m1_s10_data;    
input           m1_s11_cmd_cur; 
input           m1_s11_cmd_last; 
input           m1_s11_data;    
input           m1_s1_cmd_cur;  
input           m1_s1_cmd_last; 
input           m1_s1_data;     
input           m1_s2_cmd_cur;  
input           m1_s2_cmd_last; 
input           m1_s2_data;     
input           m1_s3_cmd_cur;  
input           m1_s3_cmd_last; 
input           m1_s3_data;     
input           m1_s4_cmd_cur;  
input           m1_s4_cmd_last; 
input           m1_s4_data;     
input           m1_s5_cmd_cur;  
input           m1_s5_cmd_last; 
input           m1_s5_data;     
input           m1_s6_cmd_cur;  
input           m1_s6_cmd_last; 
input           m1_s6_data;     
input           m1_s7_cmd_cur;  
input           m1_s7_cmd_last; 
input           m1_s7_data;     
input           m1_s8_cmd_cur;  
input           m1_s8_cmd_last; 
input           m1_s8_data;     
input           m1_s9_cmd_cur;  
input           m1_s9_cmd_last; 
input           m1_s9_data;     
input   [31:0]  m2_haddr;       
input   [2 :0]  m2_hburst;      
input   [3 :0]  m2_hprot;       
input   [2 :0]  m2_hsize;       
input   [1 :0]  m2_htrans;      
input   [31:0]  m2_hwdata;      
input           m2_hwrite;      
input           m2_latch_cmd;   
input           m2_nor_hready;  
input           m2_s0_cmd_cur;  
input           m2_s0_cmd_last; 
input           m2_s0_data;     
input           m2_s10_cmd_cur; 
input           m2_s10_cmd_last; 
input           m2_s10_data;    
input           m2_s11_cmd_cur; 
input           m2_s11_cmd_last; 
input           m2_s11_data;    
input           m2_s1_cmd_cur;  
input           m2_s1_cmd_last; 
input           m2_s1_data;     
input           m2_s2_cmd_cur;  
input           m2_s2_cmd_last; 
input           m2_s2_data;     
input           m2_s3_cmd_cur;  
input           m2_s3_cmd_last; 
input           m2_s3_data;     
input           m2_s4_cmd_cur;  
input           m2_s4_cmd_last; 
input           m2_s4_data;     
input           m2_s5_cmd_cur;  
input           m2_s5_cmd_last; 
input           m2_s5_data;     
input           m2_s6_cmd_cur;  
input           m2_s6_cmd_last; 
input           m2_s6_data;     
input           m2_s7_cmd_cur;  
input           m2_s7_cmd_last; 
input           m2_s7_data;     
input           m2_s8_cmd_cur;  
input           m2_s8_cmd_last; 
input           m2_s8_data;     
input           m2_s9_cmd_cur;  
input           m2_s9_cmd_last; 
input           m2_s9_data;     
input   [31:0]  m3_haddr;       
input   [2 :0]  m3_hburst;      
input   [3 :0]  m3_hprot;       
input   [2 :0]  m3_hsize;       
input   [1 :0]  m3_htrans;      
input   [31:0]  m3_hwdata;      
input           m3_hwrite;      
input           m3_latch_cmd;   
input           m3_nor_hready;  
input           m3_s0_cmd_cur;  
input           m3_s0_cmd_last; 
input           m3_s0_data;     
input           m3_s10_cmd_cur; 
input           m3_s10_cmd_last; 
input           m3_s10_data;    
input           m3_s11_cmd_cur; 
input           m3_s11_cmd_last; 
input           m3_s11_data;    
input           m3_s1_cmd_cur;  
input           m3_s1_cmd_last; 
input           m3_s1_data;     
input           m3_s2_cmd_cur;  
input           m3_s2_cmd_last; 
input           m3_s2_data;     
input           m3_s3_cmd_cur;  
input           m3_s3_cmd_last; 
input           m3_s3_data;     
input           m3_s4_cmd_cur;  
input           m3_s4_cmd_last; 
input           m3_s4_data;     
input           m3_s5_cmd_cur;  
input           m3_s5_cmd_last; 
input           m3_s5_data;     
input           m3_s6_cmd_cur;  
input           m3_s6_cmd_last; 
input           m3_s6_data;     
input           m3_s7_cmd_cur;  
input           m3_s7_cmd_last; 
input           m3_s7_data;     
input           m3_s8_cmd_cur;  
input           m3_s8_cmd_last; 
input           m3_s8_data;     
input           m3_s9_cmd_cur;  
input           m3_s9_cmd_last; 
input           m3_s9_data;     
input   [31:0]  m4_haddr;       
input   [2 :0]  m4_hburst;      
input   [3 :0]  m4_hprot;       
input   [2 :0]  m4_hsize;       
input   [1 :0]  m4_htrans;      
input   [31:0]  m4_hwdata;      
input           m4_hwrite;      
input           m4_latch_cmd;   
input           m4_nor_hready;  
input           m4_s0_cmd_cur;  
input           m4_s0_cmd_last; 
input           m4_s0_data;     
input           m4_s10_cmd_cur; 
input           m4_s10_cmd_last; 
input           m4_s10_data;    
input           m4_s11_cmd_cur; 
input           m4_s11_cmd_last; 
input           m4_s11_data;    
input           m4_s1_cmd_cur;  
input           m4_s1_cmd_last; 
input           m4_s1_data;     
input           m4_s2_cmd_cur;  
input           m4_s2_cmd_last; 
input           m4_s2_data;     
input           m4_s3_cmd_cur;  
input           m4_s3_cmd_last; 
input           m4_s3_data;     
input           m4_s4_cmd_cur;  
input           m4_s4_cmd_last; 
input           m4_s4_data;     
input           m4_s5_cmd_cur;  
input           m4_s5_cmd_last; 
input           m4_s5_data;     
input           m4_s6_cmd_cur;  
input           m4_s6_cmd_last; 
input           m4_s6_data;     
input           m4_s7_cmd_cur;  
input           m4_s7_cmd_last; 
input           m4_s7_data;     
input           m4_s8_cmd_cur;  
input           m4_s8_cmd_last; 
input           m4_s8_data;     
input           m4_s9_cmd_cur;  
input           m4_s9_cmd_last; 
input           m4_s9_data;     
input   [31:0]  m5_haddr;       
input   [2 :0]  m5_hburst;      
input   [3 :0]  m5_hprot;       
input   [2 :0]  m5_hsize;       
input   [1 :0]  m5_htrans;      
input   [31:0]  m5_hwdata;      
input           m5_hwrite;      
input           m5_latch_cmd;   
input           m5_nor_hready;  
input           m5_s0_cmd_cur;  
input           m5_s0_cmd_last; 
input           m5_s0_data;     
input           m5_s10_cmd_cur; 
input           m5_s10_cmd_last; 
input           m5_s10_data;    
input           m5_s11_cmd_cur; 
input           m5_s11_cmd_last; 
input           m5_s11_data;    
input           m5_s1_cmd_cur;  
input           m5_s1_cmd_last; 
input           m5_s1_data;     
input           m5_s2_cmd_cur;  
input           m5_s2_cmd_last; 
input           m5_s2_data;     
input           m5_s3_cmd_cur;  
input           m5_s3_cmd_last; 
input           m5_s3_data;     
input           m5_s4_cmd_cur;  
input           m5_s4_cmd_last; 
input           m5_s4_data;     
input           m5_s5_cmd_cur;  
input           m5_s5_cmd_last; 
input           m5_s5_data;     
input           m5_s6_cmd_cur;  
input           m5_s6_cmd_last; 
input           m5_s6_data;     
input           m5_s7_cmd_cur;  
input           m5_s7_cmd_last; 
input           m5_s7_data;     
input           m5_s8_cmd_cur;  
input           m5_s8_cmd_last; 
input           m5_s8_data;     
input           m5_s9_cmd_cur;  
input           m5_s9_cmd_last; 
input           m5_s9_data;     
input   [31:0]  m6_haddr;       
input   [2 :0]  m6_hburst;      
input   [3 :0]  m6_hprot;       
input   [2 :0]  m6_hsize;       
input   [1 :0]  m6_htrans;      
input   [31:0]  m6_hwdata;      
input           m6_hwrite;      
input           m6_latch_cmd;   
input           m6_nor_hready;  
input           m6_s0_cmd_cur;  
input           m6_s0_cmd_last; 
input           m6_s0_data;     
input           m6_s10_cmd_cur; 
input           m6_s10_cmd_last; 
input           m6_s10_data;    
input           m6_s11_cmd_cur; 
input           m6_s11_cmd_last; 
input           m6_s11_data;    
input           m6_s1_cmd_cur;  
input           m6_s1_cmd_last; 
input           m6_s1_data;     
input           m6_s2_cmd_cur;  
input           m6_s2_cmd_last; 
input           m6_s2_data;     
input           m6_s3_cmd_cur;  
input           m6_s3_cmd_last; 
input           m6_s3_data;     
input           m6_s4_cmd_cur;  
input           m6_s4_cmd_last; 
input           m6_s4_data;     
input           m6_s5_cmd_cur;  
input           m6_s5_cmd_last; 
input           m6_s5_data;     
input           m6_s6_cmd_cur;  
input           m6_s6_cmd_last; 
input           m6_s6_data;     
input           m6_s7_cmd_cur;  
input           m6_s7_cmd_last; 
input           m6_s7_data;     
input           m6_s8_cmd_cur;  
input           m6_s8_cmd_last; 
input           m6_s8_data;     
input           m6_s9_cmd_cur;  
input           m6_s9_cmd_last; 
input           m6_s9_data;     
input   [31:0]  s0_hrdata;      
input   [1 :0]  s0_hresp;       
input   [31:0]  s10_hrdata;     
input   [1 :0]  s10_hresp;      
input   [31:0]  s11_hrdata;     
input   [1 :0]  s11_hresp;      
input   [31:0]  s1_hrdata;      
input   [1 :0]  s1_hresp;       
input   [31:0]  s2_hrdata;      
input   [1 :0]  s2_hresp;       
input   [31:0]  s3_hrdata;      
input   [1 :0]  s3_hresp;       
input   [31:0]  s4_hrdata;      
input   [1 :0]  s4_hresp;       
input   [31:0]  s5_hrdata;      
input   [1 :0]  s5_hresp;       
input   [31:0]  s6_hrdata;      
input   [1 :0]  s6_hresp;       
input   [31:0]  s7_hrdata;      
input   [1 :0]  s7_hresp;       
input   [31:0]  s8_hrdata;      
input   [1 :0]  s8_hresp;       
input   [31:0]  s9_hrdata;      
input   [1 :0]  s9_hresp;       
output          m0_hgrant;      
output  [31:0]  m0_hrdata;      
output          m0_hready;      
output  [1 :0]  m0_hresp;       
output          m0_s0_req;      
output          m0_s10_req;     
output          m0_s11_req;     
output          m0_s1_req;      
output          m0_s2_req;      
output          m0_s3_req;      
output          m0_s4_req;      
output          m0_s5_req;      
output          m0_s6_req;      
output          m0_s7_req;      
output          m0_s8_req;      
output          m0_s9_req;      
output          m1_hgrant;      
output  [31:0]  m1_hrdata;      
output          m1_hready;      
output  [1 :0]  m1_hresp;       
output          m1_s0_req;      
output          m1_s10_req;     
output          m1_s11_req;     
output          m1_s1_req;      
output          m1_s2_req;      
output          m1_s3_req;      
output          m1_s4_req;      
output          m1_s5_req;      
output          m1_s6_req;      
output          m1_s7_req;      
output          m1_s8_req;      
output          m1_s9_req;      
output          m2_hgrant;      
output  [31:0]  m2_hrdata;      
output          m2_hready;      
output  [1 :0]  m2_hresp;       
output          m2_s0_req;      
output          m2_s10_req;     
output          m2_s11_req;     
output          m2_s1_req;      
output          m2_s2_req;      
output          m2_s3_req;      
output          m2_s4_req;      
output          m2_s5_req;      
output          m2_s6_req;      
output          m2_s7_req;      
output          m2_s8_req;      
output          m2_s9_req;      
output          m3_hgrant;      
output  [31:0]  m3_hrdata;      
output          m3_hready;      
output  [1 :0]  m3_hresp;       
output          m3_s0_req;      
output          m3_s10_req;     
output          m3_s11_req;     
output          m3_s1_req;      
output          m3_s2_req;      
output          m3_s3_req;      
output          m3_s4_req;      
output          m3_s5_req;      
output          m3_s6_req;      
output          m3_s7_req;      
output          m3_s8_req;      
output          m3_s9_req;      
output          m4_hgrant;      
output  [31:0]  m4_hrdata;      
output          m4_hready;      
output  [1 :0]  m4_hresp;       
output          m4_s0_req;      
output          m4_s10_req;     
output          m4_s11_req;     
output          m4_s1_req;      
output          m4_s2_req;      
output          m4_s3_req;      
output          m4_s4_req;      
output          m4_s5_req;      
output          m4_s6_req;      
output          m4_s7_req;      
output          m4_s8_req;      
output          m4_s9_req;      
output          m5_hgrant;      
output  [31:0]  m5_hrdata;      
output          m5_hready;      
output  [1 :0]  m5_hresp;       
output          m5_s0_req;      
output          m5_s10_req;     
output          m5_s11_req;     
output          m5_s1_req;      
output          m5_s2_req;      
output          m5_s3_req;      
output          m5_s4_req;      
output          m5_s5_req;      
output          m5_s6_req;      
output          m5_s7_req;      
output          m5_s8_req;      
output          m5_s9_req;      
output          m6_hgrant;      
output  [31:0]  m6_hrdata;      
output          m6_hready;      
output  [1 :0]  m6_hresp;       
output          m6_s0_req;      
output          m6_s10_req;     
output          m6_s11_req;     
output          m6_s1_req;      
output          m6_s2_req;      
output          m6_s3_req;      
output          m6_s4_req;      
output          m6_s5_req;      
output          m6_s6_req;      
output          m6_s7_req;      
output          m6_s8_req;      
output          m6_s9_req;      
output  [31:0]  s0_haddr;       
output  [2 :0]  s0_hburst;      
output  [3 :0]  s0_hprot;       
output          s0_hselx;       
output  [2 :0]  s0_hsize;       
output  [1 :0]  s0_htrans;      
output  [31:0]  s0_hwdata;      
output          s0_hwrite;      
output  [6 :0]  s0_req;         
output  [31:0]  s10_haddr;      
output  [2 :0]  s10_hburst;     
output  [3 :0]  s10_hprot;      
output          s10_hselx;      
output  [2 :0]  s10_hsize;      
output  [1 :0]  s10_htrans;     
output  [31:0]  s10_hwdata;     
output          s10_hwrite;     
output  [6 :0]  s10_req;        
output  [31:0]  s11_haddr;      
output  [2 :0]  s11_hburst;     
output  [3 :0]  s11_hprot;      
output          s11_hselx;      
output  [2 :0]  s11_hsize;      
output  [1 :0]  s11_htrans;     
output  [31:0]  s11_hwdata;     
output          s11_hwrite;     
output  [6 :0]  s11_req;        
output  [31:0]  s1_haddr;       
output  [2 :0]  s1_hburst;      
output  [3 :0]  s1_hprot;       
output          s1_hselx;       
output  [2 :0]  s1_hsize;       
output  [1 :0]  s1_htrans;      
output  [31:0]  s1_hwdata;      
output          s1_hwrite;      
output  [6 :0]  s1_req;         
output  [31:0]  s2_haddr;       
output  [2 :0]  s2_hburst;      
output  [3 :0]  s2_hprot;       
output          s2_hselx;       
output  [2 :0]  s2_hsize;       
output  [1 :0]  s2_htrans;      
output  [31:0]  s2_hwdata;      
output          s2_hwrite;      
output  [6 :0]  s2_req;         
output  [31:0]  s3_haddr;       
output  [2 :0]  s3_hburst;      
output  [3 :0]  s3_hprot;       
output          s3_hselx;       
output  [2 :0]  s3_hsize;       
output  [1 :0]  s3_htrans;      
output  [31:0]  s3_hwdata;      
output          s3_hwrite;      
output  [6 :0]  s3_req;         
output  [31:0]  s4_haddr;       
output  [2 :0]  s4_hburst;      
output  [3 :0]  s4_hprot;       
output          s4_hselx;       
output  [2 :0]  s4_hsize;       
output  [1 :0]  s4_htrans;      
output  [31:0]  s4_hwdata;      
output          s4_hwrite;      
output  [6 :0]  s4_req;         
output  [31:0]  s5_haddr;       
output  [2 :0]  s5_hburst;      
output  [3 :0]  s5_hprot;       
output          s5_hselx;       
output  [2 :0]  s5_hsize;       
output  [1 :0]  s5_htrans;      
output  [31:0]  s5_hwdata;      
output          s5_hwrite;      
output  [6 :0]  s5_req;         
output  [31:0]  s6_haddr;       
output  [2 :0]  s6_hburst;      
output  [3 :0]  s6_hprot;       
output          s6_hselx;       
output  [2 :0]  s6_hsize;       
output  [1 :0]  s6_htrans;      
output  [31:0]  s6_hwdata;      
output          s6_hwrite;      
output  [6 :0]  s6_req;         
output  [31:0]  s7_haddr;       
output  [2 :0]  s7_hburst;      
output  [3 :0]  s7_hprot;       
output          s7_hselx;       
output  [2 :0]  s7_hsize;       
output  [1 :0]  s7_htrans;      
output  [31:0]  s7_hwdata;      
output          s7_hwrite;      
output  [6 :0]  s7_req;         
output  [31:0]  s8_haddr;       
output  [2 :0]  s8_hburst;      
output  [3 :0]  s8_hprot;       
output          s8_hselx;       
output  [2 :0]  s8_hsize;       
output  [1 :0]  s8_htrans;      
output  [31:0]  s8_hwdata;      
output          s8_hwrite;      
output  [6 :0]  s8_req;         
output  [31:0]  s9_haddr;       
output  [2 :0]  s9_hburst;      
output  [3 :0]  s9_hprot;       
output          s9_hselx;       
output  [2 :0]  s9_hsize;       
output  [1 :0]  s9_htrans;      
output  [31:0]  s9_hwdata;      
output          s9_hwrite;      
output  [6 :0]  s9_req;         
reg             m0_addr_err_d;  
reg             m0_addr_err_d2; 
reg     [44:0]  m0_ctrl_bus_ff; 
reg             m1_addr_err_d;  
reg             m1_addr_err_d2; 
reg     [44:0]  m1_ctrl_bus_ff; 
reg             m2_addr_err_d;  
reg             m2_addr_err_d2; 
reg     [44:0]  m2_ctrl_bus_ff; 
reg             m3_addr_err_d;  
reg             m3_addr_err_d2; 
reg     [44:0]  m3_ctrl_bus_ff; 
reg             m4_addr_err_d;  
reg             m4_addr_err_d2; 
reg     [44:0]  m4_ctrl_bus_ff; 
reg             m5_addr_err_d;  
reg             m5_addr_err_d2; 
reg     [44:0]  m5_ctrl_bus_ff; 
reg             m6_addr_err_d;  
reg             m6_addr_err_d2; 
reg     [44:0]  m6_ctrl_bus_ff; 
wire            hclk;           
wire            hresetn;        
wire            m0_addr_err;    
wire    [44:0]  m0_ctrl_bus;    
wire            m0_err_hready;  
wire    [1 :0]  m0_err_hresp;   
wire    [31:0]  m0_haddr;       
wire    [2 :0]  m0_hburst;      
wire            m0_hgrant;      
wire    [3 :0]  m0_hprot;       
wire    [31:0]  m0_hrdata;      
wire            m0_hready;      
wire    [1 :0]  m0_hresp;       
wire    [2 :0]  m0_hsize;       
wire    [1 :0]  m0_htrans;      
wire    [31:0]  m0_hwdata;      
wire            m0_hwrite;      
wire            m0_latch_cmd;   
wire            m0_nor_hready;  
wire            m0_s0_cmd_cur;  
wire            m0_s0_cmd_last; 
wire    [44:0]  m0_s0_ctrl_bus; 
wire            m0_s0_data;     
wire            m0_s0_req;      
wire            m0_s10_cmd_cur; 
wire            m0_s10_cmd_last; 
wire    [44:0]  m0_s10_ctrl_bus; 
wire            m0_s10_data;    
wire            m0_s10_req;     
wire            m0_s11_cmd_cur; 
wire            m0_s11_cmd_last; 
wire    [44:0]  m0_s11_ctrl_bus; 
wire            m0_s11_data;    
wire            m0_s11_req;     
wire            m0_s1_cmd_cur;  
wire            m0_s1_cmd_last; 
wire    [44:0]  m0_s1_ctrl_bus; 
wire            m0_s1_data;     
wire            m0_s1_req;      
wire            m0_s2_cmd_cur;  
wire            m0_s2_cmd_last; 
wire    [44:0]  m0_s2_ctrl_bus; 
wire            m0_s2_data;     
wire            m0_s2_req;      
wire            m0_s3_cmd_cur;  
wire            m0_s3_cmd_last; 
wire    [44:0]  m0_s3_ctrl_bus; 
wire            m0_s3_data;     
wire            m0_s3_req;      
wire            m0_s4_cmd_cur;  
wire            m0_s4_cmd_last; 
wire    [44:0]  m0_s4_ctrl_bus; 
wire            m0_s4_data;     
wire            m0_s4_req;      
wire            m0_s5_cmd_cur;  
wire            m0_s5_cmd_last; 
wire    [44:0]  m0_s5_ctrl_bus; 
wire            m0_s5_data;     
wire            m0_s5_req;      
wire            m0_s6_cmd_cur;  
wire            m0_s6_cmd_last; 
wire    [44:0]  m0_s6_ctrl_bus; 
wire            m0_s6_data;     
wire            m0_s6_req;      
wire            m0_s7_cmd_cur;  
wire            m0_s7_cmd_last; 
wire    [44:0]  m0_s7_ctrl_bus; 
wire            m0_s7_data;     
wire            m0_s7_req;      
wire            m0_s8_cmd_cur;  
wire            m0_s8_cmd_last; 
wire    [44:0]  m0_s8_ctrl_bus; 
wire            m0_s8_data;     
wire            m0_s8_req;      
wire            m0_s9_cmd_cur;  
wire            m0_s9_cmd_last; 
wire    [44:0]  m0_s9_ctrl_bus; 
wire            m0_s9_data;     
wire            m0_s9_req;      
wire            m0_s_req;       
wire            m1_addr_err;    
wire    [44:0]  m1_ctrl_bus;    
wire            m1_err_hready;  
wire    [1 :0]  m1_err_hresp;   
wire    [31:0]  m1_haddr;       
wire    [2 :0]  m1_hburst;      
wire            m1_hgrant;      
wire    [3 :0]  m1_hprot;       
wire    [31:0]  m1_hrdata;      
wire            m1_hready;      
wire    [1 :0]  m1_hresp;       
wire    [2 :0]  m1_hsize;       
wire    [1 :0]  m1_htrans;      
wire    [31:0]  m1_hwdata;      
wire            m1_hwrite;      
wire            m1_latch_cmd;   
wire            m1_nor_hready;  
wire            m1_s0_cmd_cur;  
wire            m1_s0_cmd_last; 
wire    [44:0]  m1_s0_ctrl_bus; 
wire            m1_s0_data;     
wire            m1_s0_req;      
wire            m1_s10_cmd_cur; 
wire            m1_s10_cmd_last; 
wire    [44:0]  m1_s10_ctrl_bus; 
wire            m1_s10_data;    
wire            m1_s10_req;     
wire            m1_s11_cmd_cur; 
wire            m1_s11_cmd_last; 
wire    [44:0]  m1_s11_ctrl_bus; 
wire            m1_s11_data;    
wire            m1_s11_req;     
wire            m1_s1_cmd_cur;  
wire            m1_s1_cmd_last; 
wire    [44:0]  m1_s1_ctrl_bus; 
wire            m1_s1_data;     
wire            m1_s1_req;      
wire            m1_s2_cmd_cur;  
wire            m1_s2_cmd_last; 
wire    [44:0]  m1_s2_ctrl_bus; 
wire            m1_s2_data;     
wire            m1_s2_req;      
wire            m1_s3_cmd_cur;  
wire            m1_s3_cmd_last; 
wire    [44:0]  m1_s3_ctrl_bus; 
wire            m1_s3_data;     
wire            m1_s3_req;      
wire            m1_s4_cmd_cur;  
wire            m1_s4_cmd_last; 
wire    [44:0]  m1_s4_ctrl_bus; 
wire            m1_s4_data;     
wire            m1_s4_req;      
wire            m1_s5_cmd_cur;  
wire            m1_s5_cmd_last; 
wire    [44:0]  m1_s5_ctrl_bus; 
wire            m1_s5_data;     
wire            m1_s5_req;      
wire            m1_s6_cmd_cur;  
wire            m1_s6_cmd_last; 
wire    [44:0]  m1_s6_ctrl_bus; 
wire            m1_s6_data;     
wire            m1_s6_req;      
wire            m1_s7_cmd_cur;  
wire            m1_s7_cmd_last; 
wire    [44:0]  m1_s7_ctrl_bus; 
wire            m1_s7_data;     
wire            m1_s7_req;      
wire            m1_s8_cmd_cur;  
wire            m1_s8_cmd_last; 
wire    [44:0]  m1_s8_ctrl_bus; 
wire            m1_s8_data;     
wire            m1_s8_req;      
wire            m1_s9_cmd_cur;  
wire            m1_s9_cmd_last; 
wire    [44:0]  m1_s9_ctrl_bus; 
wire            m1_s9_data;     
wire            m1_s9_req;      
wire            m1_s_req;       
wire            m2_addr_err;    
wire    [44:0]  m2_ctrl_bus;    
wire            m2_err_hready;  
wire    [1 :0]  m2_err_hresp;   
wire    [31:0]  m2_haddr;       
wire    [2 :0]  m2_hburst;      
wire            m2_hgrant;      
wire    [3 :0]  m2_hprot;       
wire    [31:0]  m2_hrdata;      
wire            m2_hready;      
wire    [1 :0]  m2_hresp;       
wire    [2 :0]  m2_hsize;       
wire    [1 :0]  m2_htrans;      
wire    [31:0]  m2_hwdata;      
wire            m2_hwrite;      
wire            m2_latch_cmd;   
wire            m2_nor_hready;  
wire            m2_s0_cmd_cur;  
wire            m2_s0_cmd_last; 
wire    [44:0]  m2_s0_ctrl_bus; 
wire            m2_s0_data;     
wire            m2_s0_req;      
wire            m2_s10_cmd_cur; 
wire            m2_s10_cmd_last; 
wire    [44:0]  m2_s10_ctrl_bus; 
wire            m2_s10_data;    
wire            m2_s10_req;     
wire            m2_s11_cmd_cur; 
wire            m2_s11_cmd_last; 
wire    [44:0]  m2_s11_ctrl_bus; 
wire            m2_s11_data;    
wire            m2_s11_req;     
wire            m2_s1_cmd_cur;  
wire            m2_s1_cmd_last; 
wire    [44:0]  m2_s1_ctrl_bus; 
wire            m2_s1_data;     
wire            m2_s1_req;      
wire            m2_s2_cmd_cur;  
wire            m2_s2_cmd_last; 
wire    [44:0]  m2_s2_ctrl_bus; 
wire            m2_s2_data;     
wire            m2_s2_req;      
wire            m2_s3_cmd_cur;  
wire            m2_s3_cmd_last; 
wire    [44:0]  m2_s3_ctrl_bus; 
wire            m2_s3_data;     
wire            m2_s3_req;      
wire            m2_s4_cmd_cur;  
wire            m2_s4_cmd_last; 
wire    [44:0]  m2_s4_ctrl_bus; 
wire            m2_s4_data;     
wire            m2_s4_req;      
wire            m2_s5_cmd_cur;  
wire            m2_s5_cmd_last; 
wire    [44:0]  m2_s5_ctrl_bus; 
wire            m2_s5_data;     
wire            m2_s5_req;      
wire            m2_s6_cmd_cur;  
wire            m2_s6_cmd_last; 
wire    [44:0]  m2_s6_ctrl_bus; 
wire            m2_s6_data;     
wire            m2_s6_req;      
wire            m2_s7_cmd_cur;  
wire            m2_s7_cmd_last; 
wire    [44:0]  m2_s7_ctrl_bus; 
wire            m2_s7_data;     
wire            m2_s7_req;      
wire            m2_s8_cmd_cur;  
wire            m2_s8_cmd_last; 
wire    [44:0]  m2_s8_ctrl_bus; 
wire            m2_s8_data;     
wire            m2_s8_req;      
wire            m2_s9_cmd_cur;  
wire            m2_s9_cmd_last; 
wire    [44:0]  m2_s9_ctrl_bus; 
wire            m2_s9_data;     
wire            m2_s9_req;      
wire            m2_s_req;       
wire            m3_addr_err;    
wire    [44:0]  m3_ctrl_bus;    
wire            m3_err_hready;  
wire    [1 :0]  m3_err_hresp;   
wire    [31:0]  m3_haddr;       
wire    [2 :0]  m3_hburst;      
wire            m3_hgrant;      
wire    [3 :0]  m3_hprot;       
wire    [31:0]  m3_hrdata;      
wire            m3_hready;      
wire    [1 :0]  m3_hresp;       
wire    [2 :0]  m3_hsize;       
wire    [1 :0]  m3_htrans;      
wire    [31:0]  m3_hwdata;      
wire            m3_hwrite;      
wire            m3_latch_cmd;   
wire            m3_nor_hready;  
wire            m3_s0_cmd_cur;  
wire            m3_s0_cmd_last; 
wire    [44:0]  m3_s0_ctrl_bus; 
wire            m3_s0_data;     
wire            m3_s0_req;      
wire            m3_s10_cmd_cur; 
wire            m3_s10_cmd_last; 
wire    [44:0]  m3_s10_ctrl_bus; 
wire            m3_s10_data;    
wire            m3_s10_req;     
wire            m3_s11_cmd_cur; 
wire            m3_s11_cmd_last; 
wire    [44:0]  m3_s11_ctrl_bus; 
wire            m3_s11_data;    
wire            m3_s11_req;     
wire            m3_s1_cmd_cur;  
wire            m3_s1_cmd_last; 
wire    [44:0]  m3_s1_ctrl_bus; 
wire            m3_s1_data;     
wire            m3_s1_req;      
wire            m3_s2_cmd_cur;  
wire            m3_s2_cmd_last; 
wire    [44:0]  m3_s2_ctrl_bus; 
wire            m3_s2_data;     
wire            m3_s2_req;      
wire            m3_s3_cmd_cur;  
wire            m3_s3_cmd_last; 
wire    [44:0]  m3_s3_ctrl_bus; 
wire            m3_s3_data;     
wire            m3_s3_req;      
wire            m3_s4_cmd_cur;  
wire            m3_s4_cmd_last; 
wire    [44:0]  m3_s4_ctrl_bus; 
wire            m3_s4_data;     
wire            m3_s4_req;      
wire            m3_s5_cmd_cur;  
wire            m3_s5_cmd_last; 
wire    [44:0]  m3_s5_ctrl_bus; 
wire            m3_s5_data;     
wire            m3_s5_req;      
wire            m3_s6_cmd_cur;  
wire            m3_s6_cmd_last; 
wire    [44:0]  m3_s6_ctrl_bus; 
wire            m3_s6_data;     
wire            m3_s6_req;      
wire            m3_s7_cmd_cur;  
wire            m3_s7_cmd_last; 
wire    [44:0]  m3_s7_ctrl_bus; 
wire            m3_s7_data;     
wire            m3_s7_req;      
wire            m3_s8_cmd_cur;  
wire            m3_s8_cmd_last; 
wire    [44:0]  m3_s8_ctrl_bus; 
wire            m3_s8_data;     
wire            m3_s8_req;      
wire            m3_s9_cmd_cur;  
wire            m3_s9_cmd_last; 
wire    [44:0]  m3_s9_ctrl_bus; 
wire            m3_s9_data;     
wire            m3_s9_req;      
wire            m3_s_req;       
wire            m4_addr_err;    
wire    [44:0]  m4_ctrl_bus;    
wire            m4_err_hready;  
wire    [1 :0]  m4_err_hresp;   
wire    [31:0]  m4_haddr;       
wire    [2 :0]  m4_hburst;      
wire            m4_hgrant;      
wire    [3 :0]  m4_hprot;       
wire    [31:0]  m4_hrdata;      
wire            m4_hready;      
wire    [1 :0]  m4_hresp;       
wire    [2 :0]  m4_hsize;       
wire    [1 :0]  m4_htrans;      
wire    [31:0]  m4_hwdata;      
wire            m4_hwrite;      
wire            m4_latch_cmd;   
wire            m4_nor_hready;  
wire            m4_s0_cmd_cur;  
wire            m4_s0_cmd_last; 
wire    [44:0]  m4_s0_ctrl_bus; 
wire            m4_s0_data;     
wire            m4_s0_req;      
wire            m4_s10_cmd_cur; 
wire            m4_s10_cmd_last; 
wire    [44:0]  m4_s10_ctrl_bus; 
wire            m4_s10_data;    
wire            m4_s10_req;     
wire            m4_s11_cmd_cur; 
wire            m4_s11_cmd_last; 
wire    [44:0]  m4_s11_ctrl_bus; 
wire            m4_s11_data;    
wire            m4_s11_req;     
wire            m4_s1_cmd_cur;  
wire            m4_s1_cmd_last; 
wire    [44:0]  m4_s1_ctrl_bus; 
wire            m4_s1_data;     
wire            m4_s1_req;      
wire            m4_s2_cmd_cur;  
wire            m4_s2_cmd_last; 
wire    [44:0]  m4_s2_ctrl_bus; 
wire            m4_s2_data;     
wire            m4_s2_req;      
wire            m4_s3_cmd_cur;  
wire            m4_s3_cmd_last; 
wire    [44:0]  m4_s3_ctrl_bus; 
wire            m4_s3_data;     
wire            m4_s3_req;      
wire            m4_s4_cmd_cur;  
wire            m4_s4_cmd_last; 
wire    [44:0]  m4_s4_ctrl_bus; 
wire            m4_s4_data;     
wire            m4_s4_req;      
wire            m4_s5_cmd_cur;  
wire            m4_s5_cmd_last; 
wire    [44:0]  m4_s5_ctrl_bus; 
wire            m4_s5_data;     
wire            m4_s5_req;      
wire            m4_s6_cmd_cur;  
wire            m4_s6_cmd_last; 
wire    [44:0]  m4_s6_ctrl_bus; 
wire            m4_s6_data;     
wire            m4_s6_req;      
wire            m4_s7_cmd_cur;  
wire            m4_s7_cmd_last; 
wire    [44:0]  m4_s7_ctrl_bus; 
wire            m4_s7_data;     
wire            m4_s7_req;      
wire            m4_s8_cmd_cur;  
wire            m4_s8_cmd_last; 
wire    [44:0]  m4_s8_ctrl_bus; 
wire            m4_s8_data;     
wire            m4_s8_req;      
wire            m4_s9_cmd_cur;  
wire            m4_s9_cmd_last; 
wire    [44:0]  m4_s9_ctrl_bus; 
wire            m4_s9_data;     
wire            m4_s9_req;      
wire            m4_s_req;       
wire            m5_addr_err;    
wire    [44:0]  m5_ctrl_bus;    
wire            m5_err_hready;  
wire    [1 :0]  m5_err_hresp;   
wire    [31:0]  m5_haddr;       
wire    [2 :0]  m5_hburst;      
wire            m5_hgrant;      
wire    [3 :0]  m5_hprot;       
wire    [31:0]  m5_hrdata;      
wire            m5_hready;      
wire    [1 :0]  m5_hresp;       
wire    [2 :0]  m5_hsize;       
wire    [1 :0]  m5_htrans;      
wire    [31:0]  m5_hwdata;      
wire            m5_hwrite;      
wire            m5_latch_cmd;   
wire            m5_nor_hready;  
wire            m5_s0_cmd_cur;  
wire            m5_s0_cmd_last; 
wire    [44:0]  m5_s0_ctrl_bus; 
wire            m5_s0_data;     
wire            m5_s0_req;      
wire            m5_s10_cmd_cur; 
wire            m5_s10_cmd_last; 
wire    [44:0]  m5_s10_ctrl_bus; 
wire            m5_s10_data;    
wire            m5_s10_req;     
wire            m5_s11_cmd_cur; 
wire            m5_s11_cmd_last; 
wire    [44:0]  m5_s11_ctrl_bus; 
wire            m5_s11_data;    
wire            m5_s11_req;     
wire            m5_s1_cmd_cur;  
wire            m5_s1_cmd_last; 
wire    [44:0]  m5_s1_ctrl_bus; 
wire            m5_s1_data;     
wire            m5_s1_req;      
wire            m5_s2_cmd_cur;  
wire            m5_s2_cmd_last; 
wire    [44:0]  m5_s2_ctrl_bus; 
wire            m5_s2_data;     
wire            m5_s2_req;      
wire            m5_s3_cmd_cur;  
wire            m5_s3_cmd_last; 
wire    [44:0]  m5_s3_ctrl_bus; 
wire            m5_s3_data;     
wire            m5_s3_req;      
wire            m5_s4_cmd_cur;  
wire            m5_s4_cmd_last; 
wire    [44:0]  m5_s4_ctrl_bus; 
wire            m5_s4_data;     
wire            m5_s4_req;      
wire            m5_s5_cmd_cur;  
wire            m5_s5_cmd_last; 
wire    [44:0]  m5_s5_ctrl_bus; 
wire            m5_s5_data;     
wire            m5_s5_req;      
wire            m5_s6_cmd_cur;  
wire            m5_s6_cmd_last; 
wire    [44:0]  m5_s6_ctrl_bus; 
wire            m5_s6_data;     
wire            m5_s6_req;      
wire            m5_s7_cmd_cur;  
wire            m5_s7_cmd_last; 
wire    [44:0]  m5_s7_ctrl_bus; 
wire            m5_s7_data;     
wire            m5_s7_req;      
wire            m5_s8_cmd_cur;  
wire            m5_s8_cmd_last; 
wire    [44:0]  m5_s8_ctrl_bus; 
wire            m5_s8_data;     
wire            m5_s8_req;      
wire            m5_s9_cmd_cur;  
wire            m5_s9_cmd_last; 
wire    [44:0]  m5_s9_ctrl_bus; 
wire            m5_s9_data;     
wire            m5_s9_req;      
wire            m5_s_req;       
wire            m6_addr_err;    
wire    [44:0]  m6_ctrl_bus;    
wire            m6_err_hready;  
wire    [1 :0]  m6_err_hresp;   
wire    [31:0]  m6_haddr;       
wire    [2 :0]  m6_hburst;      
wire            m6_hgrant;      
wire    [3 :0]  m6_hprot;       
wire    [31:0]  m6_hrdata;      
wire            m6_hready;      
wire    [1 :0]  m6_hresp;       
wire    [2 :0]  m6_hsize;       
wire    [1 :0]  m6_htrans;      
wire    [31:0]  m6_hwdata;      
wire            m6_hwrite;      
wire            m6_latch_cmd;   
wire            m6_nor_hready;  
wire            m6_s0_cmd_cur;  
wire            m6_s0_cmd_last; 
wire    [44:0]  m6_s0_ctrl_bus; 
wire            m6_s0_data;     
wire            m6_s0_req;      
wire            m6_s10_cmd_cur; 
wire            m6_s10_cmd_last; 
wire    [44:0]  m6_s10_ctrl_bus; 
wire            m6_s10_data;    
wire            m6_s10_req;     
wire            m6_s11_cmd_cur; 
wire            m6_s11_cmd_last; 
wire    [44:0]  m6_s11_ctrl_bus; 
wire            m6_s11_data;    
wire            m6_s11_req;     
wire            m6_s1_cmd_cur;  
wire            m6_s1_cmd_last; 
wire    [44:0]  m6_s1_ctrl_bus; 
wire            m6_s1_data;     
wire            m6_s1_req;      
wire            m6_s2_cmd_cur;  
wire            m6_s2_cmd_last; 
wire    [44:0]  m6_s2_ctrl_bus; 
wire            m6_s2_data;     
wire            m6_s2_req;      
wire            m6_s3_cmd_cur;  
wire            m6_s3_cmd_last; 
wire    [44:0]  m6_s3_ctrl_bus; 
wire            m6_s3_data;     
wire            m6_s3_req;      
wire            m6_s4_cmd_cur;  
wire            m6_s4_cmd_last; 
wire    [44:0]  m6_s4_ctrl_bus; 
wire            m6_s4_data;     
wire            m6_s4_req;      
wire            m6_s5_cmd_cur;  
wire            m6_s5_cmd_last; 
wire    [44:0]  m6_s5_ctrl_bus; 
wire            m6_s5_data;     
wire            m6_s5_req;      
wire            m6_s6_cmd_cur;  
wire            m6_s6_cmd_last; 
wire    [44:0]  m6_s6_ctrl_bus; 
wire            m6_s6_data;     
wire            m6_s6_req;      
wire            m6_s7_cmd_cur;  
wire            m6_s7_cmd_last; 
wire    [44:0]  m6_s7_ctrl_bus; 
wire            m6_s7_data;     
wire            m6_s7_req;      
wire            m6_s8_cmd_cur;  
wire            m6_s8_cmd_last; 
wire    [44:0]  m6_s8_ctrl_bus; 
wire            m6_s8_data;     
wire            m6_s8_req;      
wire            m6_s9_cmd_cur;  
wire            m6_s9_cmd_last; 
wire    [44:0]  m6_s9_ctrl_bus; 
wire            m6_s9_data;     
wire            m6_s9_req;      
wire            m6_s_req;       
wire    [44:0]  s0_ctrl_bus;    
wire    [31:0]  s0_haddr;       
wire    [2 :0]  s0_hburst;      
wire    [3 :0]  s0_hprot;       
wire    [31:0]  s0_hrdata;      
wire    [1 :0]  s0_hresp;       
wire            s0_hselx;       
wire    [2 :0]  s0_hsize;       
wire    [1 :0]  s0_htrans;      
wire    [31:0]  s0_hwdata;      
wire            s0_hwrite;      
wire    [6 :0]  s0_req;         
wire    [44:0]  s10_ctrl_bus;   
wire    [31:0]  s10_haddr;      
wire    [2 :0]  s10_hburst;     
wire    [3 :0]  s10_hprot;      
wire    [31:0]  s10_hrdata;     
wire    [1 :0]  s10_hresp;      
wire            s10_hselx;      
wire    [2 :0]  s10_hsize;      
wire    [1 :0]  s10_htrans;     
wire    [31:0]  s10_hwdata;     
wire            s10_hwrite;     
wire    [6 :0]  s10_req;        
wire    [44:0]  s11_ctrl_bus;   
wire    [31:0]  s11_haddr;      
wire    [2 :0]  s11_hburst;     
wire    [3 :0]  s11_hprot;      
wire    [31:0]  s11_hrdata;     
wire    [1 :0]  s11_hresp;      
wire            s11_hselx;      
wire    [2 :0]  s11_hsize;      
wire    [1 :0]  s11_htrans;     
wire    [31:0]  s11_hwdata;     
wire            s11_hwrite;     
wire    [6 :0]  s11_req;        
wire    [44:0]  s1_ctrl_bus;    
wire    [31:0]  s1_haddr;       
wire    [2 :0]  s1_hburst;      
wire    [3 :0]  s1_hprot;       
wire    [31:0]  s1_hrdata;      
wire    [1 :0]  s1_hresp;       
wire            s1_hselx;       
wire    [2 :0]  s1_hsize;       
wire    [1 :0]  s1_htrans;      
wire    [31:0]  s1_hwdata;      
wire            s1_hwrite;      
wire    [6 :0]  s1_req;         
wire    [44:0]  s2_ctrl_bus;    
wire    [31:0]  s2_haddr;       
wire    [2 :0]  s2_hburst;      
wire    [3 :0]  s2_hprot;       
wire    [31:0]  s2_hrdata;      
wire    [1 :0]  s2_hresp;       
wire            s2_hselx;       
wire    [2 :0]  s2_hsize;       
wire    [1 :0]  s2_htrans;      
wire    [31:0]  s2_hwdata;      
wire            s2_hwrite;      
wire    [6 :0]  s2_req;         
wire    [44:0]  s3_ctrl_bus;    
wire    [31:0]  s3_haddr;       
wire    [2 :0]  s3_hburst;      
wire    [3 :0]  s3_hprot;       
wire    [31:0]  s3_hrdata;      
wire    [1 :0]  s3_hresp;       
wire            s3_hselx;       
wire    [2 :0]  s3_hsize;       
wire    [1 :0]  s3_htrans;      
wire    [31:0]  s3_hwdata;      
wire            s3_hwrite;      
wire    [6 :0]  s3_req;         
wire    [44:0]  s4_ctrl_bus;    
wire    [31:0]  s4_haddr;       
wire    [2 :0]  s4_hburst;      
wire    [3 :0]  s4_hprot;       
wire    [31:0]  s4_hrdata;      
wire    [1 :0]  s4_hresp;       
wire            s4_hselx;       
wire    [2 :0]  s4_hsize;       
wire    [1 :0]  s4_htrans;      
wire    [31:0]  s4_hwdata;      
wire            s4_hwrite;      
wire    [6 :0]  s4_req;         
wire    [44:0]  s5_ctrl_bus;    
wire    [31:0]  s5_haddr;       
wire    [2 :0]  s5_hburst;      
wire    [3 :0]  s5_hprot;       
wire    [31:0]  s5_hrdata;      
wire    [1 :0]  s5_hresp;       
wire            s5_hselx;       
wire    [2 :0]  s5_hsize;       
wire    [1 :0]  s5_htrans;      
wire    [31:0]  s5_hwdata;      
wire            s5_hwrite;      
wire    [6 :0]  s5_req;         
wire    [44:0]  s6_ctrl_bus;    
wire    [31:0]  s6_haddr;       
wire    [2 :0]  s6_hburst;      
wire    [3 :0]  s6_hprot;       
wire    [31:0]  s6_hrdata;      
wire    [1 :0]  s6_hresp;       
wire            s6_hselx;       
wire    [2 :0]  s6_hsize;       
wire    [1 :0]  s6_htrans;      
wire    [31:0]  s6_hwdata;      
wire            s6_hwrite;      
wire    [6 :0]  s6_req;         
wire    [44:0]  s7_ctrl_bus;    
wire    [31:0]  s7_haddr;       
wire    [2 :0]  s7_hburst;      
wire    [3 :0]  s7_hprot;       
wire    [31:0]  s7_hrdata;      
wire    [1 :0]  s7_hresp;       
wire            s7_hselx;       
wire    [2 :0]  s7_hsize;       
wire    [1 :0]  s7_htrans;      
wire    [31:0]  s7_hwdata;      
wire            s7_hwrite;      
wire    [6 :0]  s7_req;         
wire    [44:0]  s8_ctrl_bus;    
wire    [31:0]  s8_haddr;       
wire    [2 :0]  s8_hburst;      
wire    [3 :0]  s8_hprot;       
wire    [31:0]  s8_hrdata;      
wire    [1 :0]  s8_hresp;       
wire            s8_hselx;       
wire    [2 :0]  s8_hsize;       
wire    [1 :0]  s8_htrans;      
wire    [31:0]  s8_hwdata;      
wire            s8_hwrite;      
wire    [6 :0]  s8_req;         
wire    [44:0]  s9_ctrl_bus;    
wire    [31:0]  s9_haddr;       
wire    [2 :0]  s9_hburst;      
wire    [3 :0]  s9_hprot;       
wire    [31:0]  s9_hrdata;      
wire    [1 :0]  s9_hresp;       
wire            s9_hselx;       
wire    [2 :0]  s9_hsize;       
wire    [1 :0]  s9_htrans;      
wire    [31:0]  s9_hwdata;      
wire            s9_hwrite;      
wire    [6 :0]  s9_req;         
parameter BUS_WIDTH = 45;
assign m0_s0_req =( m0_haddr[31:0] >= 32'h00000000) & (m0_haddr[31:0] <= 32'h0000ffff) & (m0_htrans[1]);
assign m0_s1_req =( m0_haddr[31:0] >= 32'h10000000) & (m0_haddr[31:0] <= 32'h1007ffff) & (m0_htrans[1]);
assign m0_s2_req =( m0_haddr[31:0] >= 32'h20000000) & (m0_haddr[31:0] <= 32'h2000ffff) & (m0_htrans[1]);
assign m0_s3_req =( m0_haddr[31:0] >= 32'h20010000) & (m0_haddr[31:0] <= 32'h2001ffff) & (m0_htrans[1]);
assign m0_s4_req =( m0_haddr[31:0] >= 32'h20020000) & (m0_haddr[31:0] <= 32'h2002ffff) & (m0_htrans[1]);
assign m0_s5_req =( m0_haddr[31:0] >= 32'h30000000) & (m0_haddr[31:0] <= 32'h3fffffff) & (m0_htrans[1]);
assign m0_s6_req =( m0_haddr[31:0] >= 32'h40000000) & (m0_haddr[31:0] <= 32'h40003fff) & (m0_htrans[1]);
assign m0_s7_req =( m0_haddr[31:0] >= 32'h40010000) & (m0_haddr[31:0] <= 32'h4001ffff) & (m0_htrans[1]);
assign m0_s8_req =( m0_haddr[31:0] >= 32'h40020000) & (m0_haddr[31:0] <= 32'h4002ffff) & (m0_htrans[1]);
assign m0_s9_req =( m0_haddr[31:0] >= 32'h40100000) & (m0_haddr[31:0] <= 32'h401fffff) & (m0_htrans[1]);
assign m0_s10_req =( m0_haddr[31:0] >= 32'h40200000) & (m0_haddr[31:0] <= 32'h7fffffff) & (m0_htrans[1]);
assign m0_s11_req =( m0_haddr[31:0] >= 32'h80000000) & (m0_haddr[31:0] <= 32'h9fffffff) & (m0_htrans[1]);
assign m1_s0_req =( m1_haddr[31:0] >= 32'h00000000) & (m1_haddr[31:0] <= 32'h0000ffff) & (m1_htrans[1]);
assign m1_s1_req =( m1_haddr[31:0] >= 32'h10000000) & (m1_haddr[31:0] <= 32'h1007ffff) & (m1_htrans[1]);
assign m1_s2_req =( m1_haddr[31:0] >= 32'h20000000) & (m1_haddr[31:0] <= 32'h2000ffff) & (m1_htrans[1]);
assign m1_s3_req =( m1_haddr[31:0] >= 32'h20010000) & (m1_haddr[31:0] <= 32'h2001ffff) & (m1_htrans[1]);
assign m1_s4_req =( m1_haddr[31:0] >= 32'h20020000) & (m1_haddr[31:0] <= 32'h2002ffff) & (m1_htrans[1]);
assign m1_s5_req =( m1_haddr[31:0] >= 32'h30000000) & (m1_haddr[31:0] <= 32'h3fffffff) & (m1_htrans[1]);
assign m1_s6_req =( m1_haddr[31:0] >= 32'h40000000) & (m1_haddr[31:0] <= 32'h40003fff) & (m1_htrans[1]);
assign m1_s7_req =( m1_haddr[31:0] >= 32'h40010000) & (m1_haddr[31:0] <= 32'h4001ffff) & (m1_htrans[1]);
assign m1_s8_req =( m1_haddr[31:0] >= 32'h40020000) & (m1_haddr[31:0] <= 32'h4002ffff) & (m1_htrans[1]);
assign m1_s9_req =( m1_haddr[31:0] >= 32'h40100000) & (m1_haddr[31:0] <= 32'h401fffff) & (m1_htrans[1]);
assign m1_s10_req =( m1_haddr[31:0] >= 32'h40200000) & (m1_haddr[31:0] <= 32'h7fffffff) & (m1_htrans[1]);
assign m1_s11_req =( m1_haddr[31:0] >= 32'h80000000) & (m1_haddr[31:0] <= 32'h9fffffff) & (m1_htrans[1]);
assign m2_s0_req =( m2_haddr[31:0] >= 32'h00000000) & (m2_haddr[31:0] <= 32'h0000ffff) & (m2_htrans[1]);
assign m2_s1_req =( m2_haddr[31:0] >= 32'h10000000) & (m2_haddr[31:0] <= 32'h1007ffff) & (m2_htrans[1]);
assign m2_s2_req =( m2_haddr[31:0] >= 32'h20000000) & (m2_haddr[31:0] <= 32'h2000ffff) & (m2_htrans[1]);
assign m2_s3_req =( m2_haddr[31:0] >= 32'h20010000) & (m2_haddr[31:0] <= 32'h2001ffff) & (m2_htrans[1]);
assign m2_s4_req =( m2_haddr[31:0] >= 32'h20020000) & (m2_haddr[31:0] <= 32'h2002ffff) & (m2_htrans[1]);
assign m2_s5_req =( m2_haddr[31:0] >= 32'h30000000) & (m2_haddr[31:0] <= 32'h3fffffff) & (m2_htrans[1]);
assign m2_s6_req =( m2_haddr[31:0] >= 32'h40000000) & (m2_haddr[31:0] <= 32'h40003fff) & (m2_htrans[1]);
assign m2_s7_req =( m2_haddr[31:0] >= 32'h40010000) & (m2_haddr[31:0] <= 32'h4001ffff) & (m2_htrans[1]);
assign m2_s8_req =( m2_haddr[31:0] >= 32'h40020000) & (m2_haddr[31:0] <= 32'h4002ffff) & (m2_htrans[1]);
assign m2_s9_req =( m2_haddr[31:0] >= 32'h40100000) & (m2_haddr[31:0] <= 32'h401fffff) & (m2_htrans[1]);
assign m2_s10_req =( m2_haddr[31:0] >= 32'h40200000) & (m2_haddr[31:0] <= 32'h7fffffff) & (m2_htrans[1]);
assign m2_s11_req =( m2_haddr[31:0] >= 32'h80000000) & (m2_haddr[31:0] <= 32'h9fffffff) & (m2_htrans[1]);
assign m3_s0_req =( m3_haddr[31:0] >= 32'h00000000) & (m3_haddr[31:0] <= 32'h0000ffff) & (m3_htrans[1]);
assign m3_s1_req =( m3_haddr[31:0] >= 32'h10000000) & (m3_haddr[31:0] <= 32'h1007ffff) & (m3_htrans[1]);
assign m3_s2_req =( m3_haddr[31:0] >= 32'h20000000) & (m3_haddr[31:0] <= 32'h2000ffff) & (m3_htrans[1]);
assign m3_s3_req =( m3_haddr[31:0] >= 32'h20010000) & (m3_haddr[31:0] <= 32'h2001ffff) & (m3_htrans[1]);
assign m3_s4_req =( m3_haddr[31:0] >= 32'h20020000) & (m3_haddr[31:0] <= 32'h2002ffff) & (m3_htrans[1]);
assign m3_s5_req =( m3_haddr[31:0] >= 32'h30000000) & (m3_haddr[31:0] <= 32'h3fffffff) & (m3_htrans[1]);
assign m3_s6_req =( m3_haddr[31:0] >= 32'h40000000) & (m3_haddr[31:0] <= 32'h40003fff) & (m3_htrans[1]);
assign m3_s7_req =( m3_haddr[31:0] >= 32'h40010000) & (m3_haddr[31:0] <= 32'h4001ffff) & (m3_htrans[1]);
assign m3_s8_req =( m3_haddr[31:0] >= 32'h40020000) & (m3_haddr[31:0] <= 32'h4002ffff) & (m3_htrans[1]);
assign m3_s9_req =( m3_haddr[31:0] >= 32'h40100000) & (m3_haddr[31:0] <= 32'h401fffff) & (m3_htrans[1]);
assign m3_s10_req =( m3_haddr[31:0] >= 32'h40200000) & (m3_haddr[31:0] <= 32'h7fffffff) & (m3_htrans[1]);
assign m3_s11_req =( m3_haddr[31:0] >= 32'h80000000) & (m3_haddr[31:0] <= 32'h9fffffff) & (m3_htrans[1]);
assign m4_s0_req =( m4_haddr[31:0] >= 32'h00000000) & (m4_haddr[31:0] <= 32'h0000ffff) & (m4_htrans[1]);
assign m4_s1_req =( m4_haddr[31:0] >= 32'h10000000) & (m4_haddr[31:0] <= 32'h1007ffff) & (m4_htrans[1]);
assign m4_s2_req =( m4_haddr[31:0] >= 32'h20000000) & (m4_haddr[31:0] <= 32'h2000ffff) & (m4_htrans[1]);
assign m4_s3_req =( m4_haddr[31:0] >= 32'h20010000) & (m4_haddr[31:0] <= 32'h2001ffff) & (m4_htrans[1]);
assign m4_s4_req =( m4_haddr[31:0] >= 32'h20020000) & (m4_haddr[31:0] <= 32'h2002ffff) & (m4_htrans[1]);
assign m4_s5_req =( m4_haddr[31:0] >= 32'h30000000) & (m4_haddr[31:0] <= 32'h3fffffff) & (m4_htrans[1]);
assign m4_s6_req =( m4_haddr[31:0] >= 32'h40000000) & (m4_haddr[31:0] <= 32'h40003fff) & (m4_htrans[1]);
assign m4_s7_req =( m4_haddr[31:0] >= 32'h40010000) & (m4_haddr[31:0] <= 32'h4001ffff) & (m4_htrans[1]);
assign m4_s8_req =( m4_haddr[31:0] >= 32'h40020000) & (m4_haddr[31:0] <= 32'h4002ffff) & (m4_htrans[1]);
assign m4_s9_req =( m4_haddr[31:0] >= 32'h40100000) & (m4_haddr[31:0] <= 32'h401fffff) & (m4_htrans[1]);
assign m4_s10_req =( m4_haddr[31:0] >= 32'h40200000) & (m4_haddr[31:0] <= 32'h7fffffff) & (m4_htrans[1]);
assign m4_s11_req =( m4_haddr[31:0] >= 32'h80000000) & (m4_haddr[31:0] <= 32'h9fffffff) & (m4_htrans[1]);
assign m5_s0_req =( m5_haddr[31:0] >= 32'h00000000) & (m5_haddr[31:0] <= 32'h0000ffff) & (m5_htrans[1]);
assign m5_s1_req =( m5_haddr[31:0] >= 32'h10000000) & (m5_haddr[31:0] <= 32'h1007ffff) & (m5_htrans[1]);
assign m5_s2_req =( m5_haddr[31:0] >= 32'h20000000) & (m5_haddr[31:0] <= 32'h2000ffff) & (m5_htrans[1]);
assign m5_s3_req =( m5_haddr[31:0] >= 32'h20010000) & (m5_haddr[31:0] <= 32'h2001ffff) & (m5_htrans[1]);
assign m5_s4_req =( m5_haddr[31:0] >= 32'h20020000) & (m5_haddr[31:0] <= 32'h2002ffff) & (m5_htrans[1]);
assign m5_s5_req =( m5_haddr[31:0] >= 32'h30000000) & (m5_haddr[31:0] <= 32'h3fffffff) & (m5_htrans[1]);
assign m5_s6_req =( m5_haddr[31:0] >= 32'h40000000) & (m5_haddr[31:0] <= 32'h40003fff) & (m5_htrans[1]);
assign m5_s7_req =( m5_haddr[31:0] >= 32'h40010000) & (m5_haddr[31:0] <= 32'h4001ffff) & (m5_htrans[1]);
assign m5_s8_req =( m5_haddr[31:0] >= 32'h40020000) & (m5_haddr[31:0] <= 32'h4002ffff) & (m5_htrans[1]);
assign m5_s9_req =( m5_haddr[31:0] >= 32'h40100000) & (m5_haddr[31:0] <= 32'h401fffff) & (m5_htrans[1]);
assign m5_s10_req =( m5_haddr[31:0] >= 32'h40200000) & (m5_haddr[31:0] <= 32'h7fffffff) & (m5_htrans[1]);
assign m5_s11_req =( m5_haddr[31:0] >= 32'h80000000) & (m5_haddr[31:0] <= 32'h9fffffff) & (m5_htrans[1]);
assign m6_s0_req =( m6_haddr[31:0] >= 32'h00000000) & (m6_haddr[31:0] <= 32'h0000ffff) & (m6_htrans[1]);
assign m6_s1_req =( m6_haddr[31:0] >= 32'h10000000) & (m6_haddr[31:0] <= 32'h1007ffff) & (m6_htrans[1]);
assign m6_s2_req =( m6_haddr[31:0] >= 32'h20000000) & (m6_haddr[31:0] <= 32'h2000ffff) & (m6_htrans[1]);
assign m6_s3_req =( m6_haddr[31:0] >= 32'h20010000) & (m6_haddr[31:0] <= 32'h2001ffff) & (m6_htrans[1]);
assign m6_s4_req =( m6_haddr[31:0] >= 32'h20020000) & (m6_haddr[31:0] <= 32'h2002ffff) & (m6_htrans[1]);
assign m6_s5_req =( m6_haddr[31:0] >= 32'h30000000) & (m6_haddr[31:0] <= 32'h3fffffff) & (m6_htrans[1]);
assign m6_s6_req =( m6_haddr[31:0] >= 32'h40000000) & (m6_haddr[31:0] <= 32'h40003fff) & (m6_htrans[1]);
assign m6_s7_req =( m6_haddr[31:0] >= 32'h40010000) & (m6_haddr[31:0] <= 32'h4001ffff) & (m6_htrans[1]);
assign m6_s8_req =( m6_haddr[31:0] >= 32'h40020000) & (m6_haddr[31:0] <= 32'h4002ffff) & (m6_htrans[1]);
assign m6_s9_req =( m6_haddr[31:0] >= 32'h40100000) & (m6_haddr[31:0] <= 32'h401fffff) & (m6_htrans[1]);
assign m6_s10_req =( m6_haddr[31:0] >= 32'h40200000) & (m6_haddr[31:0] <= 32'h7fffffff) & (m6_htrans[1]);
assign m6_s11_req =( m6_haddr[31:0] >= 32'h80000000) & (m6_haddr[31:0] <= 32'h9fffffff) & (m6_htrans[1]);
assign m0_s_req = 
                    m0_s0_req |
                    m0_s1_req |
                    m0_s2_req |
                    m0_s3_req |
                    m0_s4_req |
                    m0_s5_req |
                    m0_s6_req |
                    m0_s7_req |
                    m0_s8_req |
                    m0_s9_req |
                    m0_s10_req |
                    m0_s11_req ;
assign m0_addr_err = m0_htrans[1] & (~m0_s_req) & m0_hready ;
always @ (posedge hclk or negedge hresetn)
   begin
      if(!hresetn) begin
         m0_addr_err_d <= 1'b0;
         m0_addr_err_d2 <= 1'b0;
      end
      else begin
         m0_addr_err_d <= m0_addr_err;
         m0_addr_err_d2 <= m0_addr_err_d;
      end
   end
assign m0_err_hresp[1:0] = (m0_addr_err_d|m0_addr_err_d2) ? 2'b01: 2'b00;
assign m0_err_hready = (m0_addr_err_d & (~m0_addr_err_d2));
assign m1_s_req = 
                    m1_s0_req |
                    m1_s1_req |
                    m1_s2_req |
                    m1_s3_req |
                    m1_s4_req |
                    m1_s5_req |
                    m1_s6_req |
                    m1_s7_req |
                    m1_s8_req |
                    m1_s9_req |
                    m1_s10_req |
                    m1_s11_req ;
assign m1_addr_err = m1_htrans[1] & (~m1_s_req) & m1_hready ;
always @ (posedge hclk or negedge hresetn)
   begin
      if(!hresetn) begin
         m1_addr_err_d <= 1'b0;
         m1_addr_err_d2 <= 1'b0;
      end
      else begin
         m1_addr_err_d <= m1_addr_err;
         m1_addr_err_d2 <= m1_addr_err_d;
      end
   end
assign m1_err_hresp[1:0] = (m1_addr_err_d|m1_addr_err_d2) ? 2'b01: 2'b00;
assign m1_err_hready = (m1_addr_err_d & (~m1_addr_err_d2));
assign m2_s_req = 
                    m2_s0_req |
                    m2_s1_req |
                    m2_s2_req |
                    m2_s3_req |
                    m2_s4_req |
                    m2_s5_req |
                    m2_s6_req |
                    m2_s7_req |
                    m2_s8_req |
                    m2_s9_req |
                    m2_s10_req |
                    m2_s11_req ;
assign m2_addr_err = m2_htrans[1] & (~m2_s_req) & m2_hready ;
always @ (posedge hclk or negedge hresetn)
   begin
      if(!hresetn) begin
         m2_addr_err_d <= 1'b0;
         m2_addr_err_d2 <= 1'b0;
      end
      else begin
         m2_addr_err_d <= m2_addr_err;
         m2_addr_err_d2 <= m2_addr_err_d;
      end
   end
assign m2_err_hresp[1:0] = (m2_addr_err_d|m2_addr_err_d2) ? 2'b01: 2'b00;
assign m2_err_hready = (m2_addr_err_d & (~m2_addr_err_d2));
assign m3_s_req = 
                    m3_s0_req |
                    m3_s1_req |
                    m3_s2_req |
                    m3_s3_req |
                    m3_s4_req |
                    m3_s5_req |
                    m3_s6_req |
                    m3_s7_req |
                    m3_s8_req |
                    m3_s9_req |
                    m3_s10_req |
                    m3_s11_req ;
assign m3_addr_err = m3_htrans[1] & (~m3_s_req) & m3_hready ;
always @ (posedge hclk or negedge hresetn)
   begin
      if(!hresetn) begin
         m3_addr_err_d <= 1'b0;
         m3_addr_err_d2 <= 1'b0;
      end
      else begin
         m3_addr_err_d <= m3_addr_err;
         m3_addr_err_d2 <= m3_addr_err_d;
      end
   end
assign m3_err_hresp[1:0] = (m3_addr_err_d|m3_addr_err_d2) ? 2'b01: 2'b00;
assign m3_err_hready = (m3_addr_err_d & (~m3_addr_err_d2));
assign m4_s_req = 
                    m4_s0_req |
                    m4_s1_req |
                    m4_s2_req |
                    m4_s3_req |
                    m4_s4_req |
                    m4_s5_req |
                    m4_s6_req |
                    m4_s7_req |
                    m4_s8_req |
                    m4_s9_req |
                    m4_s10_req |
                    m4_s11_req ;
assign m4_addr_err = m4_htrans[1] & (~m4_s_req) & m4_hready ;
always @ (posedge hclk or negedge hresetn)
   begin
      if(!hresetn) begin
         m4_addr_err_d <= 1'b0;
         m4_addr_err_d2 <= 1'b0;
      end
      else begin
         m4_addr_err_d <= m4_addr_err;
         m4_addr_err_d2 <= m4_addr_err_d;
      end
   end
assign m4_err_hresp[1:0] = (m4_addr_err_d|m4_addr_err_d2) ? 2'b01: 2'b00;
assign m4_err_hready = (m4_addr_err_d & (~m4_addr_err_d2));
assign m5_s_req = 
                    m5_s0_req |
                    m5_s1_req |
                    m5_s2_req |
                    m5_s3_req |
                    m5_s4_req |
                    m5_s5_req |
                    m5_s6_req |
                    m5_s7_req |
                    m5_s8_req |
                    m5_s9_req |
                    m5_s10_req |
                    m5_s11_req ;
assign m5_addr_err = m5_htrans[1] & (~m5_s_req) & m5_hready ;
always @ (posedge hclk or negedge hresetn)
   begin
      if(!hresetn) begin
         m5_addr_err_d <= 1'b0;
         m5_addr_err_d2 <= 1'b0;
      end
      else begin
         m5_addr_err_d <= m5_addr_err;
         m5_addr_err_d2 <= m5_addr_err_d;
      end
   end
assign m5_err_hresp[1:0] = (m5_addr_err_d|m5_addr_err_d2) ? 2'b01: 2'b00;
assign m5_err_hready = (m5_addr_err_d & (~m5_addr_err_d2));
assign m6_s_req = 
                    m6_s0_req |
                    m6_s1_req |
                    m6_s2_req |
                    m6_s3_req |
                    m6_s4_req |
                    m6_s5_req |
                    m6_s6_req |
                    m6_s7_req |
                    m6_s8_req |
                    m6_s9_req |
                    m6_s10_req |
                    m6_s11_req ;
assign m6_addr_err = m6_htrans[1] & (~m6_s_req) & m6_hready ;
always @ (posedge hclk or negedge hresetn)
   begin
      if(!hresetn) begin
         m6_addr_err_d <= 1'b0;
         m6_addr_err_d2 <= 1'b0;
      end
      else begin
         m6_addr_err_d <= m6_addr_err;
         m6_addr_err_d2 <= m6_addr_err_d;
      end
   end
assign m6_err_hresp[1:0] = (m6_addr_err_d|m6_addr_err_d2) ? 2'b01: 2'b00;
assign m6_err_hready = (m6_addr_err_d & (~m6_addr_err_d2));
assign s0_req[7-1:0] = {
                        m0_s0_req,
                        m1_s0_req,
                        m2_s0_req,
                        m3_s0_req,
                        m4_s0_req,
                        m5_s0_req,
                        m6_s0_req};
assign s1_req[7-1:0] = {
                        m0_s1_req,
                        m1_s1_req,
                        m2_s1_req,
                        m3_s1_req,
                        m4_s1_req,
                        m5_s1_req,
                        m6_s1_req};
assign s2_req[7-1:0] = {
                        m0_s2_req,
                        m1_s2_req,
                        m2_s2_req,
                        m3_s2_req,
                        m4_s2_req,
                        m5_s2_req,
                        m6_s2_req};
assign s3_req[7-1:0] = {
                        m0_s3_req,
                        m1_s3_req,
                        m2_s3_req,
                        m3_s3_req,
                        m4_s3_req,
                        m5_s3_req,
                        m6_s3_req};
assign s4_req[7-1:0] = {
                        m0_s4_req,
                        m1_s4_req,
                        m2_s4_req,
                        m3_s4_req,
                        m4_s4_req,
                        m5_s4_req,
                        m6_s4_req};
assign s5_req[7-1:0] = {
                        m0_s5_req,
                        m1_s5_req,
                        m2_s5_req,
                        m3_s5_req,
                        m4_s5_req,
                        m5_s5_req,
                        m6_s5_req};
assign s6_req[7-1:0] = {
                        m0_s6_req,
                        m1_s6_req,
                        m2_s6_req,
                        m3_s6_req,
                        m4_s6_req,
                        m5_s6_req,
                        m6_s6_req};
assign s7_req[7-1:0] = {
                        m0_s7_req,
                        m1_s7_req,
                        m2_s7_req,
                        m3_s7_req,
                        m4_s7_req,
                        m5_s7_req,
                        m6_s7_req};
assign s8_req[7-1:0] = {
                        m0_s8_req,
                        m1_s8_req,
                        m2_s8_req,
                        m3_s8_req,
                        m4_s8_req,
                        m5_s8_req,
                        m6_s8_req};
assign s9_req[7-1:0] = {
                        m0_s9_req,
                        m1_s9_req,
                        m2_s9_req,
                        m3_s9_req,
                        m4_s9_req,
                        m5_s9_req,
                        m6_s9_req};
assign s10_req[7-1:0] = {
                        m0_s10_req,
                        m1_s10_req,
                        m2_s10_req,
                        m3_s10_req,
                        m4_s10_req,
                        m5_s10_req,
                        m6_s10_req};
assign s11_req[7-1:0] = {
                        m0_s11_req,
                        m1_s11_req,
                        m2_s11_req,
                        m3_s11_req,
                        m4_s11_req,
                        m5_s11_req,
                        m6_s11_req};
assign m0_ctrl_bus[BUS_WIDTH-1:0] = {m0_haddr[32-1:0],m0_htrans[1:0],m0_hsize[2:0],m0_hburst[2:0],m0_hprot[3:0],m0_hwrite};
assign m1_ctrl_bus[BUS_WIDTH-1:0] = {m1_haddr[32-1:0],m1_htrans[1:0],m1_hsize[2:0],m1_hburst[2:0],m1_hprot[3:0],m1_hwrite};
assign m2_ctrl_bus[BUS_WIDTH-1:0] = {m2_haddr[32-1:0],m2_htrans[1:0],m2_hsize[2:0],m2_hburst[2:0],m2_hprot[3:0],m2_hwrite};
assign m3_ctrl_bus[BUS_WIDTH-1:0] = {m3_haddr[32-1:0],m3_htrans[1:0],m3_hsize[2:0],m3_hburst[2:0],m3_hprot[3:0],m3_hwrite};
assign m4_ctrl_bus[BUS_WIDTH-1:0] = {m4_haddr[32-1:0],m4_htrans[1:0],m4_hsize[2:0],m4_hburst[2:0],m4_hprot[3:0],m4_hwrite};
assign m5_ctrl_bus[BUS_WIDTH-1:0] = {m5_haddr[32-1:0],m5_htrans[1:0],m5_hsize[2:0],m5_hburst[2:0],m5_hprot[3:0],m5_hwrite};
assign m6_ctrl_bus[BUS_WIDTH-1:0] = {m6_haddr[32-1:0],m6_htrans[1:0],m6_hsize[2:0],m6_hburst[2:0],m6_hprot[3:0],m6_hwrite};
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
       m0_ctrl_bus_ff[BUS_WIDTH-1:0] <= 0;
    else if(m0_latch_cmd)
       m0_ctrl_bus_ff[BUS_WIDTH-1:0] <= m0_ctrl_bus[BUS_WIDTH-1:0];
  end
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
       m1_ctrl_bus_ff[BUS_WIDTH-1:0] <= 0;
    else if(m1_latch_cmd)
       m1_ctrl_bus_ff[BUS_WIDTH-1:0] <= m1_ctrl_bus[BUS_WIDTH-1:0];
  end
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
       m2_ctrl_bus_ff[BUS_WIDTH-1:0] <= 0;
    else if(m2_latch_cmd)
       m2_ctrl_bus_ff[BUS_WIDTH-1:0] <= m2_ctrl_bus[BUS_WIDTH-1:0];
  end
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
       m3_ctrl_bus_ff[BUS_WIDTH-1:0] <= 0;
    else if(m3_latch_cmd)
       m3_ctrl_bus_ff[BUS_WIDTH-1:0] <= m3_ctrl_bus[BUS_WIDTH-1:0];
  end
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
       m4_ctrl_bus_ff[BUS_WIDTH-1:0] <= 0;
    else if(m4_latch_cmd)
       m4_ctrl_bus_ff[BUS_WIDTH-1:0] <= m4_ctrl_bus[BUS_WIDTH-1:0];
  end
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
       m5_ctrl_bus_ff[BUS_WIDTH-1:0] <= 0;
    else if(m5_latch_cmd)
       m5_ctrl_bus_ff[BUS_WIDTH-1:0] <= m5_ctrl_bus[BUS_WIDTH-1:0];
  end
always @ (posedge hclk or negedge hresetn)
  begin
    if(!hresetn)
       m6_ctrl_bus_ff[BUS_WIDTH-1:0] <= 0;
    else if(m6_latch_cmd)
       m6_ctrl_bus_ff[BUS_WIDTH-1:0] <= m6_ctrl_bus[BUS_WIDTH-1:0];
  end
assign m0_s0_ctrl_bus[BUS_WIDTH-1:0] = m0_s0_cmd_cur  ?  m0_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m0_s0_cmd_last ?  m0_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m0_s1_ctrl_bus[BUS_WIDTH-1:0] = m0_s1_cmd_cur  ?  m0_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m0_s1_cmd_last ?  m0_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m0_s2_ctrl_bus[BUS_WIDTH-1:0] = m0_s2_cmd_cur  ?  m0_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m0_s2_cmd_last ?  m0_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m0_s3_ctrl_bus[BUS_WIDTH-1:0] = m0_s3_cmd_cur  ?  m0_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m0_s3_cmd_last ?  m0_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m0_s4_ctrl_bus[BUS_WIDTH-1:0] = m0_s4_cmd_cur  ?  m0_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m0_s4_cmd_last ?  m0_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m0_s5_ctrl_bus[BUS_WIDTH-1:0] = m0_s5_cmd_cur  ?  m0_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m0_s5_cmd_last ?  m0_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m0_s6_ctrl_bus[BUS_WIDTH-1:0] = m0_s6_cmd_cur  ?  m0_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m0_s6_cmd_last ?  m0_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m0_s7_ctrl_bus[BUS_WIDTH-1:0] = m0_s7_cmd_cur  ?  m0_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m0_s7_cmd_last ?  m0_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m0_s8_ctrl_bus[BUS_WIDTH-1:0] = m0_s8_cmd_cur  ?  m0_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m0_s8_cmd_last ?  m0_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m0_s9_ctrl_bus[BUS_WIDTH-1:0] = m0_s9_cmd_cur  ?  m0_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m0_s9_cmd_last ?  m0_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m0_s10_ctrl_bus[BUS_WIDTH-1:0] = m0_s10_cmd_cur  ?  m0_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m0_s10_cmd_last ?  m0_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m0_s11_ctrl_bus[BUS_WIDTH-1:0] = m0_s11_cmd_cur  ?  m0_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m0_s11_cmd_last ?  m0_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m1_s0_ctrl_bus[BUS_WIDTH-1:0] = m1_s0_cmd_cur  ?  m1_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m1_s0_cmd_last ?  m1_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m1_s1_ctrl_bus[BUS_WIDTH-1:0] = m1_s1_cmd_cur  ?  m1_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m1_s1_cmd_last ?  m1_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m1_s2_ctrl_bus[BUS_WIDTH-1:0] = m1_s2_cmd_cur  ?  m1_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m1_s2_cmd_last ?  m1_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m1_s3_ctrl_bus[BUS_WIDTH-1:0] = m1_s3_cmd_cur  ?  m1_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m1_s3_cmd_last ?  m1_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m1_s4_ctrl_bus[BUS_WIDTH-1:0] = m1_s4_cmd_cur  ?  m1_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m1_s4_cmd_last ?  m1_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m1_s5_ctrl_bus[BUS_WIDTH-1:0] = m1_s5_cmd_cur  ?  m1_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m1_s5_cmd_last ?  m1_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m1_s6_ctrl_bus[BUS_WIDTH-1:0] = m1_s6_cmd_cur  ?  m1_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m1_s6_cmd_last ?  m1_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m1_s7_ctrl_bus[BUS_WIDTH-1:0] = m1_s7_cmd_cur  ?  m1_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m1_s7_cmd_last ?  m1_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m1_s8_ctrl_bus[BUS_WIDTH-1:0] = m1_s8_cmd_cur  ?  m1_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m1_s8_cmd_last ?  m1_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m1_s9_ctrl_bus[BUS_WIDTH-1:0] = m1_s9_cmd_cur  ?  m1_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m1_s9_cmd_last ?  m1_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m1_s10_ctrl_bus[BUS_WIDTH-1:0] = m1_s10_cmd_cur  ?  m1_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m1_s10_cmd_last ?  m1_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m1_s11_ctrl_bus[BUS_WIDTH-1:0] = m1_s11_cmd_cur  ?  m1_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m1_s11_cmd_last ?  m1_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m2_s0_ctrl_bus[BUS_WIDTH-1:0] = m2_s0_cmd_cur  ?  m2_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m2_s0_cmd_last ?  m2_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m2_s1_ctrl_bus[BUS_WIDTH-1:0] = m2_s1_cmd_cur  ?  m2_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m2_s1_cmd_last ?  m2_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m2_s2_ctrl_bus[BUS_WIDTH-1:0] = m2_s2_cmd_cur  ?  m2_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m2_s2_cmd_last ?  m2_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m2_s3_ctrl_bus[BUS_WIDTH-1:0] = m2_s3_cmd_cur  ?  m2_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m2_s3_cmd_last ?  m2_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m2_s4_ctrl_bus[BUS_WIDTH-1:0] = m2_s4_cmd_cur  ?  m2_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m2_s4_cmd_last ?  m2_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m2_s5_ctrl_bus[BUS_WIDTH-1:0] = m2_s5_cmd_cur  ?  m2_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m2_s5_cmd_last ?  m2_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m2_s6_ctrl_bus[BUS_WIDTH-1:0] = m2_s6_cmd_cur  ?  m2_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m2_s6_cmd_last ?  m2_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m2_s7_ctrl_bus[BUS_WIDTH-1:0] = m2_s7_cmd_cur  ?  m2_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m2_s7_cmd_last ?  m2_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m2_s8_ctrl_bus[BUS_WIDTH-1:0] = m2_s8_cmd_cur  ?  m2_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m2_s8_cmd_last ?  m2_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m2_s9_ctrl_bus[BUS_WIDTH-1:0] = m2_s9_cmd_cur  ?  m2_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m2_s9_cmd_last ?  m2_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m2_s10_ctrl_bus[BUS_WIDTH-1:0] = m2_s10_cmd_cur  ?  m2_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m2_s10_cmd_last ?  m2_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m2_s11_ctrl_bus[BUS_WIDTH-1:0] = m2_s11_cmd_cur  ?  m2_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m2_s11_cmd_last ?  m2_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m3_s0_ctrl_bus[BUS_WIDTH-1:0] = m3_s0_cmd_cur  ?  m3_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m3_s0_cmd_last ?  m3_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m3_s1_ctrl_bus[BUS_WIDTH-1:0] = m3_s1_cmd_cur  ?  m3_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m3_s1_cmd_last ?  m3_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m3_s2_ctrl_bus[BUS_WIDTH-1:0] = m3_s2_cmd_cur  ?  m3_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m3_s2_cmd_last ?  m3_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m3_s3_ctrl_bus[BUS_WIDTH-1:0] = m3_s3_cmd_cur  ?  m3_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m3_s3_cmd_last ?  m3_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m3_s4_ctrl_bus[BUS_WIDTH-1:0] = m3_s4_cmd_cur  ?  m3_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m3_s4_cmd_last ?  m3_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m3_s5_ctrl_bus[BUS_WIDTH-1:0] = m3_s5_cmd_cur  ?  m3_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m3_s5_cmd_last ?  m3_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m3_s6_ctrl_bus[BUS_WIDTH-1:0] = m3_s6_cmd_cur  ?  m3_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m3_s6_cmd_last ?  m3_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m3_s7_ctrl_bus[BUS_WIDTH-1:0] = m3_s7_cmd_cur  ?  m3_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m3_s7_cmd_last ?  m3_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m3_s8_ctrl_bus[BUS_WIDTH-1:0] = m3_s8_cmd_cur  ?  m3_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m3_s8_cmd_last ?  m3_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m3_s9_ctrl_bus[BUS_WIDTH-1:0] = m3_s9_cmd_cur  ?  m3_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m3_s9_cmd_last ?  m3_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m3_s10_ctrl_bus[BUS_WIDTH-1:0] = m3_s10_cmd_cur  ?  m3_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m3_s10_cmd_last ?  m3_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m3_s11_ctrl_bus[BUS_WIDTH-1:0] = m3_s11_cmd_cur  ?  m3_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m3_s11_cmd_last ?  m3_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m4_s0_ctrl_bus[BUS_WIDTH-1:0] = m4_s0_cmd_cur  ?  m4_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m4_s0_cmd_last ?  m4_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m4_s1_ctrl_bus[BUS_WIDTH-1:0] = m4_s1_cmd_cur  ?  m4_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m4_s1_cmd_last ?  m4_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m4_s2_ctrl_bus[BUS_WIDTH-1:0] = m4_s2_cmd_cur  ?  m4_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m4_s2_cmd_last ?  m4_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m4_s3_ctrl_bus[BUS_WIDTH-1:0] = m4_s3_cmd_cur  ?  m4_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m4_s3_cmd_last ?  m4_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m4_s4_ctrl_bus[BUS_WIDTH-1:0] = m4_s4_cmd_cur  ?  m4_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m4_s4_cmd_last ?  m4_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m4_s5_ctrl_bus[BUS_WIDTH-1:0] = m4_s5_cmd_cur  ?  m4_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m4_s5_cmd_last ?  m4_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m4_s6_ctrl_bus[BUS_WIDTH-1:0] = m4_s6_cmd_cur  ?  m4_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m4_s6_cmd_last ?  m4_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m4_s7_ctrl_bus[BUS_WIDTH-1:0] = m4_s7_cmd_cur  ?  m4_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m4_s7_cmd_last ?  m4_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m4_s8_ctrl_bus[BUS_WIDTH-1:0] = m4_s8_cmd_cur  ?  m4_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m4_s8_cmd_last ?  m4_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m4_s9_ctrl_bus[BUS_WIDTH-1:0] = m4_s9_cmd_cur  ?  m4_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m4_s9_cmd_last ?  m4_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m4_s10_ctrl_bus[BUS_WIDTH-1:0] = m4_s10_cmd_cur  ?  m4_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m4_s10_cmd_last ?  m4_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m4_s11_ctrl_bus[BUS_WIDTH-1:0] = m4_s11_cmd_cur  ?  m4_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m4_s11_cmd_last ?  m4_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m5_s0_ctrl_bus[BUS_WIDTH-1:0] = m5_s0_cmd_cur  ?  m5_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m5_s0_cmd_last ?  m5_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m5_s1_ctrl_bus[BUS_WIDTH-1:0] = m5_s1_cmd_cur  ?  m5_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m5_s1_cmd_last ?  m5_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m5_s2_ctrl_bus[BUS_WIDTH-1:0] = m5_s2_cmd_cur  ?  m5_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m5_s2_cmd_last ?  m5_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m5_s3_ctrl_bus[BUS_WIDTH-1:0] = m5_s3_cmd_cur  ?  m5_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m5_s3_cmd_last ?  m5_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m5_s4_ctrl_bus[BUS_WIDTH-1:0] = m5_s4_cmd_cur  ?  m5_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m5_s4_cmd_last ?  m5_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m5_s5_ctrl_bus[BUS_WIDTH-1:0] = m5_s5_cmd_cur  ?  m5_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m5_s5_cmd_last ?  m5_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m5_s6_ctrl_bus[BUS_WIDTH-1:0] = m5_s6_cmd_cur  ?  m5_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m5_s6_cmd_last ?  m5_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m5_s7_ctrl_bus[BUS_WIDTH-1:0] = m5_s7_cmd_cur  ?  m5_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m5_s7_cmd_last ?  m5_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m5_s8_ctrl_bus[BUS_WIDTH-1:0] = m5_s8_cmd_cur  ?  m5_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m5_s8_cmd_last ?  m5_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m5_s9_ctrl_bus[BUS_WIDTH-1:0] = m5_s9_cmd_cur  ?  m5_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m5_s9_cmd_last ?  m5_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m5_s10_ctrl_bus[BUS_WIDTH-1:0] = m5_s10_cmd_cur  ?  m5_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m5_s10_cmd_last ?  m5_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m5_s11_ctrl_bus[BUS_WIDTH-1:0] = m5_s11_cmd_cur  ?  m5_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m5_s11_cmd_last ?  m5_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m6_s0_ctrl_bus[BUS_WIDTH-1:0] = m6_s0_cmd_cur  ?  m6_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m6_s0_cmd_last ?  m6_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m6_s1_ctrl_bus[BUS_WIDTH-1:0] = m6_s1_cmd_cur  ?  m6_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m6_s1_cmd_last ?  m6_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m6_s2_ctrl_bus[BUS_WIDTH-1:0] = m6_s2_cmd_cur  ?  m6_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m6_s2_cmd_last ?  m6_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m6_s3_ctrl_bus[BUS_WIDTH-1:0] = m6_s3_cmd_cur  ?  m6_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m6_s3_cmd_last ?  m6_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m6_s4_ctrl_bus[BUS_WIDTH-1:0] = m6_s4_cmd_cur  ?  m6_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m6_s4_cmd_last ?  m6_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m6_s5_ctrl_bus[BUS_WIDTH-1:0] = m6_s5_cmd_cur  ?  m6_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m6_s5_cmd_last ?  m6_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m6_s6_ctrl_bus[BUS_WIDTH-1:0] = m6_s6_cmd_cur  ?  m6_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m6_s6_cmd_last ?  m6_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m6_s7_ctrl_bus[BUS_WIDTH-1:0] = m6_s7_cmd_cur  ?  m6_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m6_s7_cmd_last ?  m6_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m6_s8_ctrl_bus[BUS_WIDTH-1:0] = m6_s8_cmd_cur  ?  m6_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m6_s8_cmd_last ?  m6_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m6_s9_ctrl_bus[BUS_WIDTH-1:0] = m6_s9_cmd_cur  ?  m6_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m6_s9_cmd_last ?  m6_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m6_s10_ctrl_bus[BUS_WIDTH-1:0] = m6_s10_cmd_cur  ?  m6_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m6_s10_cmd_last ?  m6_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign m6_s11_ctrl_bus[BUS_WIDTH-1:0] = m6_s11_cmd_cur  ?  m6_ctrl_bus[BUS_WIDTH-1:0] : 
                                       m6_s11_cmd_last ?  m6_ctrl_bus_ff[BUS_WIDTH-1:0] : 0;
assign s0_ctrl_bus[BUS_WIDTH-1:0] = 
                                    m0_s0_ctrl_bus[BUS_WIDTH-1:0] |
                                    m1_s0_ctrl_bus[BUS_WIDTH-1:0] |
                                    m2_s0_ctrl_bus[BUS_WIDTH-1:0] |
                                    m3_s0_ctrl_bus[BUS_WIDTH-1:0] |
                                    m4_s0_ctrl_bus[BUS_WIDTH-1:0] |
                                    m5_s0_ctrl_bus[BUS_WIDTH-1:0] |
                                    m6_s0_ctrl_bus[BUS_WIDTH-1:0];
assign s1_ctrl_bus[BUS_WIDTH-1:0] = 
                                    m0_s1_ctrl_bus[BUS_WIDTH-1:0] |
                                    m1_s1_ctrl_bus[BUS_WIDTH-1:0] |
                                    m2_s1_ctrl_bus[BUS_WIDTH-1:0] |
                                    m3_s1_ctrl_bus[BUS_WIDTH-1:0] |
                                    m4_s1_ctrl_bus[BUS_WIDTH-1:0] |
                                    m5_s1_ctrl_bus[BUS_WIDTH-1:0] |
                                    m6_s1_ctrl_bus[BUS_WIDTH-1:0];
assign s2_ctrl_bus[BUS_WIDTH-1:0] = 
                                    m0_s2_ctrl_bus[BUS_WIDTH-1:0] |
                                    m1_s2_ctrl_bus[BUS_WIDTH-1:0] |
                                    m2_s2_ctrl_bus[BUS_WIDTH-1:0] |
                                    m3_s2_ctrl_bus[BUS_WIDTH-1:0] |
                                    m4_s2_ctrl_bus[BUS_WIDTH-1:0] |
                                    m5_s2_ctrl_bus[BUS_WIDTH-1:0] |
                                    m6_s2_ctrl_bus[BUS_WIDTH-1:0];
assign s3_ctrl_bus[BUS_WIDTH-1:0] = 
                                    m0_s3_ctrl_bus[BUS_WIDTH-1:0] |
                                    m1_s3_ctrl_bus[BUS_WIDTH-1:0] |
                                    m2_s3_ctrl_bus[BUS_WIDTH-1:0] |
                                    m3_s3_ctrl_bus[BUS_WIDTH-1:0] |
                                    m4_s3_ctrl_bus[BUS_WIDTH-1:0] |
                                    m5_s3_ctrl_bus[BUS_WIDTH-1:0] |
                                    m6_s3_ctrl_bus[BUS_WIDTH-1:0];
assign s4_ctrl_bus[BUS_WIDTH-1:0] = 
                                    m0_s4_ctrl_bus[BUS_WIDTH-1:0] |
                                    m1_s4_ctrl_bus[BUS_WIDTH-1:0] |
                                    m2_s4_ctrl_bus[BUS_WIDTH-1:0] |
                                    m3_s4_ctrl_bus[BUS_WIDTH-1:0] |
                                    m4_s4_ctrl_bus[BUS_WIDTH-1:0] |
                                    m5_s4_ctrl_bus[BUS_WIDTH-1:0] |
                                    m6_s4_ctrl_bus[BUS_WIDTH-1:0];
assign s5_ctrl_bus[BUS_WIDTH-1:0] = 
                                    m0_s5_ctrl_bus[BUS_WIDTH-1:0] |
                                    m1_s5_ctrl_bus[BUS_WIDTH-1:0] |
                                    m2_s5_ctrl_bus[BUS_WIDTH-1:0] |
                                    m3_s5_ctrl_bus[BUS_WIDTH-1:0] |
                                    m4_s5_ctrl_bus[BUS_WIDTH-1:0] |
                                    m5_s5_ctrl_bus[BUS_WIDTH-1:0] |
                                    m6_s5_ctrl_bus[BUS_WIDTH-1:0];
assign s6_ctrl_bus[BUS_WIDTH-1:0] = 
                                    m0_s6_ctrl_bus[BUS_WIDTH-1:0] |
                                    m1_s6_ctrl_bus[BUS_WIDTH-1:0] |
                                    m2_s6_ctrl_bus[BUS_WIDTH-1:0] |
                                    m3_s6_ctrl_bus[BUS_WIDTH-1:0] |
                                    m4_s6_ctrl_bus[BUS_WIDTH-1:0] |
                                    m5_s6_ctrl_bus[BUS_WIDTH-1:0] |
                                    m6_s6_ctrl_bus[BUS_WIDTH-1:0];
assign s7_ctrl_bus[BUS_WIDTH-1:0] = 
                                    m0_s7_ctrl_bus[BUS_WIDTH-1:0] |
                                    m1_s7_ctrl_bus[BUS_WIDTH-1:0] |
                                    m2_s7_ctrl_bus[BUS_WIDTH-1:0] |
                                    m3_s7_ctrl_bus[BUS_WIDTH-1:0] |
                                    m4_s7_ctrl_bus[BUS_WIDTH-1:0] |
                                    m5_s7_ctrl_bus[BUS_WIDTH-1:0] |
                                    m6_s7_ctrl_bus[BUS_WIDTH-1:0];
assign s8_ctrl_bus[BUS_WIDTH-1:0] = 
                                    m0_s8_ctrl_bus[BUS_WIDTH-1:0] |
                                    m1_s8_ctrl_bus[BUS_WIDTH-1:0] |
                                    m2_s8_ctrl_bus[BUS_WIDTH-1:0] |
                                    m3_s8_ctrl_bus[BUS_WIDTH-1:0] |
                                    m4_s8_ctrl_bus[BUS_WIDTH-1:0] |
                                    m5_s8_ctrl_bus[BUS_WIDTH-1:0] |
                                    m6_s8_ctrl_bus[BUS_WIDTH-1:0];
assign s9_ctrl_bus[BUS_WIDTH-1:0] = 
                                    m0_s9_ctrl_bus[BUS_WIDTH-1:0] |
                                    m1_s9_ctrl_bus[BUS_WIDTH-1:0] |
                                    m2_s9_ctrl_bus[BUS_WIDTH-1:0] |
                                    m3_s9_ctrl_bus[BUS_WIDTH-1:0] |
                                    m4_s9_ctrl_bus[BUS_WIDTH-1:0] |
                                    m5_s9_ctrl_bus[BUS_WIDTH-1:0] |
                                    m6_s9_ctrl_bus[BUS_WIDTH-1:0];
assign s10_ctrl_bus[BUS_WIDTH-1:0] = 
                                    m0_s10_ctrl_bus[BUS_WIDTH-1:0] |
                                    m1_s10_ctrl_bus[BUS_WIDTH-1:0] |
                                    m2_s10_ctrl_bus[BUS_WIDTH-1:0] |
                                    m3_s10_ctrl_bus[BUS_WIDTH-1:0] |
                                    m4_s10_ctrl_bus[BUS_WIDTH-1:0] |
                                    m5_s10_ctrl_bus[BUS_WIDTH-1:0] |
                                    m6_s10_ctrl_bus[BUS_WIDTH-1:0];
assign s11_ctrl_bus[BUS_WIDTH-1:0] = 
                                    m0_s11_ctrl_bus[BUS_WIDTH-1:0] |
                                    m1_s11_ctrl_bus[BUS_WIDTH-1:0] |
                                    m2_s11_ctrl_bus[BUS_WIDTH-1:0] |
                                    m3_s11_ctrl_bus[BUS_WIDTH-1:0] |
                                    m4_s11_ctrl_bus[BUS_WIDTH-1:0] |
                                    m5_s11_ctrl_bus[BUS_WIDTH-1:0] |
                                    m6_s11_ctrl_bus[BUS_WIDTH-1:0];
assign {s0_haddr[31:0],s0_htrans[1:0],s0_hsize[2:0],s0_hburst[2:0],s0_hprot[3:0],s0_hwrite} = s0_ctrl_bus[BUS_WIDTH-1:0];
assign {s1_haddr[31:0],s1_htrans[1:0],s1_hsize[2:0],s1_hburst[2:0],s1_hprot[3:0],s1_hwrite} = s1_ctrl_bus[BUS_WIDTH-1:0];
assign {s2_haddr[31:0],s2_htrans[1:0],s2_hsize[2:0],s2_hburst[2:0],s2_hprot[3:0],s2_hwrite} = s2_ctrl_bus[BUS_WIDTH-1:0];
assign {s3_haddr[31:0],s3_htrans[1:0],s3_hsize[2:0],s3_hburst[2:0],s3_hprot[3:0],s3_hwrite} = s3_ctrl_bus[BUS_WIDTH-1:0];
assign {s4_haddr[31:0],s4_htrans[1:0],s4_hsize[2:0],s4_hburst[2:0],s4_hprot[3:0],s4_hwrite} = s4_ctrl_bus[BUS_WIDTH-1:0];
assign {s5_haddr[31:0],s5_htrans[1:0],s5_hsize[2:0],s5_hburst[2:0],s5_hprot[3:0],s5_hwrite} = s5_ctrl_bus[BUS_WIDTH-1:0];
assign {s6_haddr[31:0],s6_htrans[1:0],s6_hsize[2:0],s6_hburst[2:0],s6_hprot[3:0],s6_hwrite} = s6_ctrl_bus[BUS_WIDTH-1:0];
assign {s7_haddr[31:0],s7_htrans[1:0],s7_hsize[2:0],s7_hburst[2:0],s7_hprot[3:0],s7_hwrite} = s7_ctrl_bus[BUS_WIDTH-1:0];
assign {s8_haddr[31:0],s8_htrans[1:0],s8_hsize[2:0],s8_hburst[2:0],s8_hprot[3:0],s8_hwrite} = s8_ctrl_bus[BUS_WIDTH-1:0];
assign {s9_haddr[31:0],s9_htrans[1:0],s9_hsize[2:0],s9_hburst[2:0],s9_hprot[3:0],s9_hwrite} = s9_ctrl_bus[BUS_WIDTH-1:0];
assign {s10_haddr[31:0],s10_htrans[1:0],s10_hsize[2:0],s10_hburst[2:0],s10_hprot[3:0],s10_hwrite} = s10_ctrl_bus[BUS_WIDTH-1:0];
assign {s11_haddr[31:0],s11_htrans[1:0],s11_hsize[2:0],s11_hburst[2:0],s11_hprot[3:0],s11_hwrite} = s11_ctrl_bus[BUS_WIDTH-1:0];
assign s0_hwdata[31:0] = 
                           (m0_hwdata[31:0] & {32{m0_s0_data}}) |
                           (m1_hwdata[31:0] & {32{m1_s0_data}}) |
                           (m2_hwdata[31:0] & {32{m2_s0_data}}) |
                           (m3_hwdata[31:0] & {32{m3_s0_data}}) |
                           (m4_hwdata[31:0] & {32{m4_s0_data}}) |
                           (m5_hwdata[31:0] & {32{m5_s0_data}}) |
                           (m6_hwdata[31:0] & {32{m6_s0_data}});
assign s1_hwdata[31:0] = 
                           (m0_hwdata[31:0] & {32{m0_s1_data}}) |
                           (m1_hwdata[31:0] & {32{m1_s1_data}}) |
                           (m2_hwdata[31:0] & {32{m2_s1_data}}) |
                           (m3_hwdata[31:0] & {32{m3_s1_data}}) |
                           (m4_hwdata[31:0] & {32{m4_s1_data}}) |
                           (m5_hwdata[31:0] & {32{m5_s1_data}}) |
                           (m6_hwdata[31:0] & {32{m6_s1_data}});
assign s2_hwdata[31:0] = 
                           (m0_hwdata[31:0] & {32{m0_s2_data}}) |
                           (m1_hwdata[31:0] & {32{m1_s2_data}}) |
                           (m2_hwdata[31:0] & {32{m2_s2_data}}) |
                           (m3_hwdata[31:0] & {32{m3_s2_data}}) |
                           (m4_hwdata[31:0] & {32{m4_s2_data}}) |
                           (m5_hwdata[31:0] & {32{m5_s2_data}}) |
                           (m6_hwdata[31:0] & {32{m6_s2_data}});
assign s3_hwdata[31:0] = 
                           (m0_hwdata[31:0] & {32{m0_s3_data}}) |
                           (m1_hwdata[31:0] & {32{m1_s3_data}}) |
                           (m2_hwdata[31:0] & {32{m2_s3_data}}) |
                           (m3_hwdata[31:0] & {32{m3_s3_data}}) |
                           (m4_hwdata[31:0] & {32{m4_s3_data}}) |
                           (m5_hwdata[31:0] & {32{m5_s3_data}}) |
                           (m6_hwdata[31:0] & {32{m6_s3_data}});
assign s4_hwdata[31:0] = 
                           (m0_hwdata[31:0] & {32{m0_s4_data}}) |
                           (m1_hwdata[31:0] & {32{m1_s4_data}}) |
                           (m2_hwdata[31:0] & {32{m2_s4_data}}) |
                           (m3_hwdata[31:0] & {32{m3_s4_data}}) |
                           (m4_hwdata[31:0] & {32{m4_s4_data}}) |
                           (m5_hwdata[31:0] & {32{m5_s4_data}}) |
                           (m6_hwdata[31:0] & {32{m6_s4_data}});
assign s5_hwdata[31:0] = 
                           (m0_hwdata[31:0] & {32{m0_s5_data}}) |
                           (m1_hwdata[31:0] & {32{m1_s5_data}}) |
                           (m2_hwdata[31:0] & {32{m2_s5_data}}) |
                           (m3_hwdata[31:0] & {32{m3_s5_data}}) |
                           (m4_hwdata[31:0] & {32{m4_s5_data}}) |
                           (m5_hwdata[31:0] & {32{m5_s5_data}}) |
                           (m6_hwdata[31:0] & {32{m6_s5_data}});
assign s6_hwdata[31:0] = 
                           (m0_hwdata[31:0] & {32{m0_s6_data}}) |
                           (m1_hwdata[31:0] & {32{m1_s6_data}}) |
                           (m2_hwdata[31:0] & {32{m2_s6_data}}) |
                           (m3_hwdata[31:0] & {32{m3_s6_data}}) |
                           (m4_hwdata[31:0] & {32{m4_s6_data}}) |
                           (m5_hwdata[31:0] & {32{m5_s6_data}}) |
                           (m6_hwdata[31:0] & {32{m6_s6_data}});
assign s7_hwdata[31:0] = 
                           (m0_hwdata[31:0] & {32{m0_s7_data}}) |
                           (m1_hwdata[31:0] & {32{m1_s7_data}}) |
                           (m2_hwdata[31:0] & {32{m2_s7_data}}) |
                           (m3_hwdata[31:0] & {32{m3_s7_data}}) |
                           (m4_hwdata[31:0] & {32{m4_s7_data}}) |
                           (m5_hwdata[31:0] & {32{m5_s7_data}}) |
                           (m6_hwdata[31:0] & {32{m6_s7_data}});
assign s8_hwdata[31:0] = 
                           (m0_hwdata[31:0] & {32{m0_s8_data}}) |
                           (m1_hwdata[31:0] & {32{m1_s8_data}}) |
                           (m2_hwdata[31:0] & {32{m2_s8_data}}) |
                           (m3_hwdata[31:0] & {32{m3_s8_data}}) |
                           (m4_hwdata[31:0] & {32{m4_s8_data}}) |
                           (m5_hwdata[31:0] & {32{m5_s8_data}}) |
                           (m6_hwdata[31:0] & {32{m6_s8_data}});
assign s9_hwdata[31:0] = 
                           (m0_hwdata[31:0] & {32{m0_s9_data}}) |
                           (m1_hwdata[31:0] & {32{m1_s9_data}}) |
                           (m2_hwdata[31:0] & {32{m2_s9_data}}) |
                           (m3_hwdata[31:0] & {32{m3_s9_data}}) |
                           (m4_hwdata[31:0] & {32{m4_s9_data}}) |
                           (m5_hwdata[31:0] & {32{m5_s9_data}}) |
                           (m6_hwdata[31:0] & {32{m6_s9_data}});
assign s10_hwdata[31:0] = 
                           (m0_hwdata[31:0] & {32{m0_s10_data}}) |
                           (m1_hwdata[31:0] & {32{m1_s10_data}}) |
                           (m2_hwdata[31:0] & {32{m2_s10_data}}) |
                           (m3_hwdata[31:0] & {32{m3_s10_data}}) |
                           (m4_hwdata[31:0] & {32{m4_s10_data}}) |
                           (m5_hwdata[31:0] & {32{m5_s10_data}}) |
                           (m6_hwdata[31:0] & {32{m6_s10_data}});
assign s11_hwdata[31:0] = 
                           (m0_hwdata[31:0] & {32{m0_s11_data}}) |
                           (m1_hwdata[31:0] & {32{m1_s11_data}}) |
                           (m2_hwdata[31:0] & {32{m2_s11_data}}) |
                           (m3_hwdata[31:0] & {32{m3_s11_data}}) |
                           (m4_hwdata[31:0] & {32{m4_s11_data}}) |
                           (m5_hwdata[31:0] & {32{m5_s11_data}}) |
                           (m6_hwdata[31:0] & {32{m6_s11_data}});
assign m0_hrdata[32-1:0] = 
                           (s0_hrdata[32-1:0] & {32{m0_s0_data}}) |
                           (s1_hrdata[32-1:0] & {32{m0_s1_data}}) |
                           (s2_hrdata[32-1:0] & {32{m0_s2_data}}) |
                           (s3_hrdata[32-1:0] & {32{m0_s3_data}}) |
                           (s4_hrdata[32-1:0] & {32{m0_s4_data}}) |
                           (s5_hrdata[32-1:0] & {32{m0_s5_data}}) |
                           (s6_hrdata[32-1:0] & {32{m0_s6_data}}) |
                           (s7_hrdata[32-1:0] & {32{m0_s7_data}}) |
                           (s8_hrdata[32-1:0] & {32{m0_s8_data}}) |
                           (s9_hrdata[32-1:0] & {32{m0_s9_data}}) |
                           (s10_hrdata[32-1:0] & {32{m0_s10_data}}) |
                           (s11_hrdata[32-1:0] & {32{m0_s11_data}});
assign m1_hrdata[32-1:0] = 
                           (s0_hrdata[32-1:0] & {32{m1_s0_data}}) |
                           (s1_hrdata[32-1:0] & {32{m1_s1_data}}) |
                           (s2_hrdata[32-1:0] & {32{m1_s2_data}}) |
                           (s3_hrdata[32-1:0] & {32{m1_s3_data}}) |
                           (s4_hrdata[32-1:0] & {32{m1_s4_data}}) |
                           (s5_hrdata[32-1:0] & {32{m1_s5_data}}) |
                           (s6_hrdata[32-1:0] & {32{m1_s6_data}}) |
                           (s7_hrdata[32-1:0] & {32{m1_s7_data}}) |
                           (s8_hrdata[32-1:0] & {32{m1_s8_data}}) |
                           (s9_hrdata[32-1:0] & {32{m1_s9_data}}) |
                           (s10_hrdata[32-1:0] & {32{m1_s10_data}}) |
                           (s11_hrdata[32-1:0] & {32{m1_s11_data}});
assign m2_hrdata[32-1:0] = 
                           (s0_hrdata[32-1:0] & {32{m2_s0_data}}) |
                           (s1_hrdata[32-1:0] & {32{m2_s1_data}}) |
                           (s2_hrdata[32-1:0] & {32{m2_s2_data}}) |
                           (s3_hrdata[32-1:0] & {32{m2_s3_data}}) |
                           (s4_hrdata[32-1:0] & {32{m2_s4_data}}) |
                           (s5_hrdata[32-1:0] & {32{m2_s5_data}}) |
                           (s6_hrdata[32-1:0] & {32{m2_s6_data}}) |
                           (s7_hrdata[32-1:0] & {32{m2_s7_data}}) |
                           (s8_hrdata[32-1:0] & {32{m2_s8_data}}) |
                           (s9_hrdata[32-1:0] & {32{m2_s9_data}}) |
                           (s10_hrdata[32-1:0] & {32{m2_s10_data}}) |
                           (s11_hrdata[32-1:0] & {32{m2_s11_data}});
assign m3_hrdata[32-1:0] = 
                           (s0_hrdata[32-1:0] & {32{m3_s0_data}}) |
                           (s1_hrdata[32-1:0] & {32{m3_s1_data}}) |
                           (s2_hrdata[32-1:0] & {32{m3_s2_data}}) |
                           (s3_hrdata[32-1:0] & {32{m3_s3_data}}) |
                           (s4_hrdata[32-1:0] & {32{m3_s4_data}}) |
                           (s5_hrdata[32-1:0] & {32{m3_s5_data}}) |
                           (s6_hrdata[32-1:0] & {32{m3_s6_data}}) |
                           (s7_hrdata[32-1:0] & {32{m3_s7_data}}) |
                           (s8_hrdata[32-1:0] & {32{m3_s8_data}}) |
                           (s9_hrdata[32-1:0] & {32{m3_s9_data}}) |
                           (s10_hrdata[32-1:0] & {32{m3_s10_data}}) |
                           (s11_hrdata[32-1:0] & {32{m3_s11_data}});
assign m4_hrdata[32-1:0] = 
                           (s0_hrdata[32-1:0] & {32{m4_s0_data}}) |
                           (s1_hrdata[32-1:0] & {32{m4_s1_data}}) |
                           (s2_hrdata[32-1:0] & {32{m4_s2_data}}) |
                           (s3_hrdata[32-1:0] & {32{m4_s3_data}}) |
                           (s4_hrdata[32-1:0] & {32{m4_s4_data}}) |
                           (s5_hrdata[32-1:0] & {32{m4_s5_data}}) |
                           (s6_hrdata[32-1:0] & {32{m4_s6_data}}) |
                           (s7_hrdata[32-1:0] & {32{m4_s7_data}}) |
                           (s8_hrdata[32-1:0] & {32{m4_s8_data}}) |
                           (s9_hrdata[32-1:0] & {32{m4_s9_data}}) |
                           (s10_hrdata[32-1:0] & {32{m4_s10_data}}) |
                           (s11_hrdata[32-1:0] & {32{m4_s11_data}});
assign m5_hrdata[32-1:0] = 
                           (s0_hrdata[32-1:0] & {32{m5_s0_data}}) |
                           (s1_hrdata[32-1:0] & {32{m5_s1_data}}) |
                           (s2_hrdata[32-1:0] & {32{m5_s2_data}}) |
                           (s3_hrdata[32-1:0] & {32{m5_s3_data}}) |
                           (s4_hrdata[32-1:0] & {32{m5_s4_data}}) |
                           (s5_hrdata[32-1:0] & {32{m5_s5_data}}) |
                           (s6_hrdata[32-1:0] & {32{m5_s6_data}}) |
                           (s7_hrdata[32-1:0] & {32{m5_s7_data}}) |
                           (s8_hrdata[32-1:0] & {32{m5_s8_data}}) |
                           (s9_hrdata[32-1:0] & {32{m5_s9_data}}) |
                           (s10_hrdata[32-1:0] & {32{m5_s10_data}}) |
                           (s11_hrdata[32-1:0] & {32{m5_s11_data}});
assign m6_hrdata[32-1:0] = 
                           (s0_hrdata[32-1:0] & {32{m6_s0_data}}) |
                           (s1_hrdata[32-1:0] & {32{m6_s1_data}}) |
                           (s2_hrdata[32-1:0] & {32{m6_s2_data}}) |
                           (s3_hrdata[32-1:0] & {32{m6_s3_data}}) |
                           (s4_hrdata[32-1:0] & {32{m6_s4_data}}) |
                           (s5_hrdata[32-1:0] & {32{m6_s5_data}}) |
                           (s6_hrdata[32-1:0] & {32{m6_s6_data}}) |
                           (s7_hrdata[32-1:0] & {32{m6_s7_data}}) |
                           (s8_hrdata[32-1:0] & {32{m6_s8_data}}) |
                           (s9_hrdata[32-1:0] & {32{m6_s9_data}}) |
                           (s10_hrdata[32-1:0] & {32{m6_s10_data}}) |
                           (s11_hrdata[32-1:0] & {32{m6_s11_data}});
assign m0_hresp[1:0] = 
                       (s0_hresp[1:0] & {2{m0_s0_data}}) |
                       (s1_hresp[1:0] & {2{m0_s1_data}}) |
                       (s2_hresp[1:0] & {2{m0_s2_data}}) |
                       (s3_hresp[1:0] & {2{m0_s3_data}}) |
                       (s4_hresp[1:0] & {2{m0_s4_data}}) |
                       (s5_hresp[1:0] & {2{m0_s5_data}}) |
                       (s6_hresp[1:0] & {2{m0_s6_data}}) |
                       (s7_hresp[1:0] & {2{m0_s7_data}}) |
                       (s8_hresp[1:0] & {2{m0_s8_data}}) |
                       (s9_hresp[1:0] & {2{m0_s9_data}}) |
                       (s10_hresp[1:0] & {2{m0_s10_data}}) |
                       (s11_hresp[1:0] & {2{m0_s11_data}}) |
                       m0_err_hresp[1:0];
assign m1_hresp[1:0] = 
                       (s0_hresp[1:0] & {2{m1_s0_data}}) |
                       (s1_hresp[1:0] & {2{m1_s1_data}}) |
                       (s2_hresp[1:0] & {2{m1_s2_data}}) |
                       (s3_hresp[1:0] & {2{m1_s3_data}}) |
                       (s4_hresp[1:0] & {2{m1_s4_data}}) |
                       (s5_hresp[1:0] & {2{m1_s5_data}}) |
                       (s6_hresp[1:0] & {2{m1_s6_data}}) |
                       (s7_hresp[1:0] & {2{m1_s7_data}}) |
                       (s8_hresp[1:0] & {2{m1_s8_data}}) |
                       (s9_hresp[1:0] & {2{m1_s9_data}}) |
                       (s10_hresp[1:0] & {2{m1_s10_data}}) |
                       (s11_hresp[1:0] & {2{m1_s11_data}}) |
                       m1_err_hresp[1:0];
assign m2_hresp[1:0] = 
                       (s0_hresp[1:0] & {2{m2_s0_data}}) |
                       (s1_hresp[1:0] & {2{m2_s1_data}}) |
                       (s2_hresp[1:0] & {2{m2_s2_data}}) |
                       (s3_hresp[1:0] & {2{m2_s3_data}}) |
                       (s4_hresp[1:0] & {2{m2_s4_data}}) |
                       (s5_hresp[1:0] & {2{m2_s5_data}}) |
                       (s6_hresp[1:0] & {2{m2_s6_data}}) |
                       (s7_hresp[1:0] & {2{m2_s7_data}}) |
                       (s8_hresp[1:0] & {2{m2_s8_data}}) |
                       (s9_hresp[1:0] & {2{m2_s9_data}}) |
                       (s10_hresp[1:0] & {2{m2_s10_data}}) |
                       (s11_hresp[1:0] & {2{m2_s11_data}}) |
                       m2_err_hresp[1:0];
assign m3_hresp[1:0] = 
                       (s0_hresp[1:0] & {2{m3_s0_data}}) |
                       (s1_hresp[1:0] & {2{m3_s1_data}}) |
                       (s2_hresp[1:0] & {2{m3_s2_data}}) |
                       (s3_hresp[1:0] & {2{m3_s3_data}}) |
                       (s4_hresp[1:0] & {2{m3_s4_data}}) |
                       (s5_hresp[1:0] & {2{m3_s5_data}}) |
                       (s6_hresp[1:0] & {2{m3_s6_data}}) |
                       (s7_hresp[1:0] & {2{m3_s7_data}}) |
                       (s8_hresp[1:0] & {2{m3_s8_data}}) |
                       (s9_hresp[1:0] & {2{m3_s9_data}}) |
                       (s10_hresp[1:0] & {2{m3_s10_data}}) |
                       (s11_hresp[1:0] & {2{m3_s11_data}}) |
                       m3_err_hresp[1:0];
assign m4_hresp[1:0] = 
                       (s0_hresp[1:0] & {2{m4_s0_data}}) |
                       (s1_hresp[1:0] & {2{m4_s1_data}}) |
                       (s2_hresp[1:0] & {2{m4_s2_data}}) |
                       (s3_hresp[1:0] & {2{m4_s3_data}}) |
                       (s4_hresp[1:0] & {2{m4_s4_data}}) |
                       (s5_hresp[1:0] & {2{m4_s5_data}}) |
                       (s6_hresp[1:0] & {2{m4_s6_data}}) |
                       (s7_hresp[1:0] & {2{m4_s7_data}}) |
                       (s8_hresp[1:0] & {2{m4_s8_data}}) |
                       (s9_hresp[1:0] & {2{m4_s9_data}}) |
                       (s10_hresp[1:0] & {2{m4_s10_data}}) |
                       (s11_hresp[1:0] & {2{m4_s11_data}}) |
                       m4_err_hresp[1:0];
assign m5_hresp[1:0] = 
                       (s0_hresp[1:0] & {2{m5_s0_data}}) |
                       (s1_hresp[1:0] & {2{m5_s1_data}}) |
                       (s2_hresp[1:0] & {2{m5_s2_data}}) |
                       (s3_hresp[1:0] & {2{m5_s3_data}}) |
                       (s4_hresp[1:0] & {2{m5_s4_data}}) |
                       (s5_hresp[1:0] & {2{m5_s5_data}}) |
                       (s6_hresp[1:0] & {2{m5_s6_data}}) |
                       (s7_hresp[1:0] & {2{m5_s7_data}}) |
                       (s8_hresp[1:0] & {2{m5_s8_data}}) |
                       (s9_hresp[1:0] & {2{m5_s9_data}}) |
                       (s10_hresp[1:0] & {2{m5_s10_data}}) |
                       (s11_hresp[1:0] & {2{m5_s11_data}}) |
                       m5_err_hresp[1:0];
assign m6_hresp[1:0] = 
                       (s0_hresp[1:0] & {2{m6_s0_data}}) |
                       (s1_hresp[1:0] & {2{m6_s1_data}}) |
                       (s2_hresp[1:0] & {2{m6_s2_data}}) |
                       (s3_hresp[1:0] & {2{m6_s3_data}}) |
                       (s4_hresp[1:0] & {2{m6_s4_data}}) |
                       (s5_hresp[1:0] & {2{m6_s5_data}}) |
                       (s6_hresp[1:0] & {2{m6_s6_data}}) |
                       (s7_hresp[1:0] & {2{m6_s7_data}}) |
                       (s8_hresp[1:0] & {2{m6_s8_data}}) |
                       (s9_hresp[1:0] & {2{m6_s9_data}}) |
                       (s10_hresp[1:0] & {2{m6_s10_data}}) |
                       (s11_hresp[1:0] & {2{m6_s11_data}}) |
                       m6_err_hresp[1:0];
assign m0_hready = (~m0_err_hready) & m0_nor_hready;
assign m1_hready = (~m1_err_hready) & m1_nor_hready;
assign m2_hready = (~m2_err_hready) & m2_nor_hready;
assign m3_hready = (~m3_err_hready) & m3_nor_hready;
assign m4_hready = (~m4_err_hready) & m4_nor_hready;
assign m5_hready = (~m5_err_hready) & m5_nor_hready;
assign m6_hready = (~m6_err_hready) & m6_nor_hready;
assign s0_hselx = 
                  m0_s0_cmd_last | m0_s0_cmd_cur |
                  m1_s0_cmd_last | m1_s0_cmd_cur |
                  m2_s0_cmd_last | m2_s0_cmd_cur |
                  m3_s0_cmd_last | m3_s0_cmd_cur |
                  m4_s0_cmd_last | m4_s0_cmd_cur |
                  m5_s0_cmd_last | m5_s0_cmd_cur |
                  m6_s0_cmd_last | m6_s0_cmd_cur;
assign s1_hselx = 
                  m0_s1_cmd_last | m0_s1_cmd_cur |
                  m1_s1_cmd_last | m1_s1_cmd_cur |
                  m2_s1_cmd_last | m2_s1_cmd_cur |
                  m3_s1_cmd_last | m3_s1_cmd_cur |
                  m4_s1_cmd_last | m4_s1_cmd_cur |
                  m5_s1_cmd_last | m5_s1_cmd_cur |
                  m6_s1_cmd_last | m6_s1_cmd_cur;
assign s2_hselx = 
                  m0_s2_cmd_last | m0_s2_cmd_cur |
                  m1_s2_cmd_last | m1_s2_cmd_cur |
                  m2_s2_cmd_last | m2_s2_cmd_cur |
                  m3_s2_cmd_last | m3_s2_cmd_cur |
                  m4_s2_cmd_last | m4_s2_cmd_cur |
                  m5_s2_cmd_last | m5_s2_cmd_cur |
                  m6_s2_cmd_last | m6_s2_cmd_cur;
assign s3_hselx = 
                  m0_s3_cmd_last | m0_s3_cmd_cur |
                  m1_s3_cmd_last | m1_s3_cmd_cur |
                  m2_s3_cmd_last | m2_s3_cmd_cur |
                  m3_s3_cmd_last | m3_s3_cmd_cur |
                  m4_s3_cmd_last | m4_s3_cmd_cur |
                  m5_s3_cmd_last | m5_s3_cmd_cur |
                  m6_s3_cmd_last | m6_s3_cmd_cur;
assign s4_hselx = 
                  m0_s4_cmd_last | m0_s4_cmd_cur |
                  m1_s4_cmd_last | m1_s4_cmd_cur |
                  m2_s4_cmd_last | m2_s4_cmd_cur |
                  m3_s4_cmd_last | m3_s4_cmd_cur |
                  m4_s4_cmd_last | m4_s4_cmd_cur |
                  m5_s4_cmd_last | m5_s4_cmd_cur |
                  m6_s4_cmd_last | m6_s4_cmd_cur;
assign s5_hselx = 
                  m0_s5_cmd_last | m0_s5_cmd_cur |
                  m1_s5_cmd_last | m1_s5_cmd_cur |
                  m2_s5_cmd_last | m2_s5_cmd_cur |
                  m3_s5_cmd_last | m3_s5_cmd_cur |
                  m4_s5_cmd_last | m4_s5_cmd_cur |
                  m5_s5_cmd_last | m5_s5_cmd_cur |
                  m6_s5_cmd_last | m6_s5_cmd_cur;
assign s6_hselx = 
                  m0_s6_cmd_last | m0_s6_cmd_cur |
                  m1_s6_cmd_last | m1_s6_cmd_cur |
                  m2_s6_cmd_last | m2_s6_cmd_cur |
                  m3_s6_cmd_last | m3_s6_cmd_cur |
                  m4_s6_cmd_last | m4_s6_cmd_cur |
                  m5_s6_cmd_last | m5_s6_cmd_cur |
                  m6_s6_cmd_last | m6_s6_cmd_cur;
assign s7_hselx = 
                  m0_s7_cmd_last | m0_s7_cmd_cur |
                  m1_s7_cmd_last | m1_s7_cmd_cur |
                  m2_s7_cmd_last | m2_s7_cmd_cur |
                  m3_s7_cmd_last | m3_s7_cmd_cur |
                  m4_s7_cmd_last | m4_s7_cmd_cur |
                  m5_s7_cmd_last | m5_s7_cmd_cur |
                  m6_s7_cmd_last | m6_s7_cmd_cur;
assign s8_hselx = 
                  m0_s8_cmd_last | m0_s8_cmd_cur |
                  m1_s8_cmd_last | m1_s8_cmd_cur |
                  m2_s8_cmd_last | m2_s8_cmd_cur |
                  m3_s8_cmd_last | m3_s8_cmd_cur |
                  m4_s8_cmd_last | m4_s8_cmd_cur |
                  m5_s8_cmd_last | m5_s8_cmd_cur |
                  m6_s8_cmd_last | m6_s8_cmd_cur;
assign s9_hselx = 
                  m0_s9_cmd_last | m0_s9_cmd_cur |
                  m1_s9_cmd_last | m1_s9_cmd_cur |
                  m2_s9_cmd_last | m2_s9_cmd_cur |
                  m3_s9_cmd_last | m3_s9_cmd_cur |
                  m4_s9_cmd_last | m4_s9_cmd_cur |
                  m5_s9_cmd_last | m5_s9_cmd_cur |
                  m6_s9_cmd_last | m6_s9_cmd_cur;
assign s10_hselx = 
                  m0_s10_cmd_last | m0_s10_cmd_cur |
                  m1_s10_cmd_last | m1_s10_cmd_cur |
                  m2_s10_cmd_last | m2_s10_cmd_cur |
                  m3_s10_cmd_last | m3_s10_cmd_cur |
                  m4_s10_cmd_last | m4_s10_cmd_cur |
                  m5_s10_cmd_last | m5_s10_cmd_cur |
                  m6_s10_cmd_last | m6_s10_cmd_cur;
assign s11_hselx = 
                  m0_s11_cmd_last | m0_s11_cmd_cur |
                  m1_s11_cmd_last | m1_s11_cmd_cur |
                  m2_s11_cmd_last | m2_s11_cmd_cur |
                  m3_s11_cmd_last | m3_s11_cmd_cur |
                  m4_s11_cmd_last | m4_s11_cmd_cur |
                  m5_s11_cmd_last | m5_s11_cmd_cur |
                  m6_s11_cmd_last | m6_s11_cmd_cur;
assign m0_hgrant = 1'b1;
assign m1_hgrant = 1'b1;
assign m2_hgrant = 1'b1;
assign m3_hgrant = 1'b1;
assign m4_hgrant = 1'b1;
assign m5_hgrant = 1'b1;
assign m6_hgrant = 1'b1;
endmodule
module ahb_matrix_7_12_main(
  hclk,
  hresetn,
  m0_haddr,
  m0_hburst,
  m0_hgrant,
  m0_hprot,
  m0_hrdata,
  m0_hready,
  m0_hresp,
  m0_hsize,
  m0_htrans,
  m0_hwdata,
  m0_hwrite,
  m1_haddr,
  m1_hburst,
  m1_hgrant,
  m1_hprot,
  m1_hrdata,
  m1_hready,
  m1_hresp,
  m1_hsize,
  m1_htrans,
  m1_hwdata,
  m1_hwrite,
  m2_haddr,
  m2_hburst,
  m2_hgrant,
  m2_hprot,
  m2_hrdata,
  m2_hready,
  m2_hresp,
  m2_hsize,
  m2_htrans,
  m2_hwdata,
  m2_hwrite,
  m3_haddr,
  m3_hburst,
  m3_hgrant,
  m3_hprot,
  m3_hrdata,
  m3_hready,
  m3_hresp,
  m3_hsize,
  m3_htrans,
  m3_hwdata,
  m3_hwrite,
  m4_haddr,
  m4_hburst,
  m4_hgrant,
  m4_hprot,
  m4_hrdata,
  m4_hready,
  m4_hresp,
  m4_hsize,
  m4_htrans,
  m4_hwdata,
  m4_hwrite,
  m5_haddr,
  m5_hburst,
  m5_hgrant,
  m5_hprot,
  m5_hrdata,
  m5_hready,
  m5_hresp,
  m5_hsize,
  m5_htrans,
  m5_hwdata,
  m5_hwrite,
  m6_haddr,
  m6_hburst,
  m6_hgrant,
  m6_hprot,
  m6_hrdata,
  m6_hready,
  m6_hresp,
  m6_hsize,
  m6_htrans,
  m6_hwdata,
  m6_hwrite,
  s0_haddr,
  s0_hburst,
  s0_hprot,
  s0_hrdata,
  s0_hready,
  s0_hresp,
  s0_hselx,
  s0_hsize,
  s0_htrans,
  s0_hwdata,
  s0_hwrite,
  s10_haddr,
  s10_hburst,
  s10_hprot,
  s10_hrdata,
  s10_hready,
  s10_hresp,
  s10_hselx,
  s10_hsize,
  s10_htrans,
  s10_hwdata,
  s10_hwrite,
  s11_haddr,
  s11_hburst,
  s11_hprot,
  s11_hrdata,
  s11_hready,
  s11_hresp,
  s11_hselx,
  s11_hsize,
  s11_htrans,
  s11_hwdata,
  s11_hwrite,
  s1_haddr,
  s1_hburst,
  s1_hprot,
  s1_hrdata,
  s1_hready,
  s1_hresp,
  s1_hselx,
  s1_hsize,
  s1_htrans,
  s1_hwdata,
  s1_hwrite,
  s2_haddr,
  s2_hburst,
  s2_hprot,
  s2_hrdata,
  s2_hready,
  s2_hresp,
  s2_hselx,
  s2_hsize,
  s2_htrans,
  s2_hwdata,
  s2_hwrite,
  s3_haddr,
  s3_hburst,
  s3_hprot,
  s3_hrdata,
  s3_hready,
  s3_hresp,
  s3_hselx,
  s3_hsize,
  s3_htrans,
  s3_hwdata,
  s3_hwrite,
  s4_haddr,
  s4_hburst,
  s4_hprot,
  s4_hrdata,
  s4_hready,
  s4_hresp,
  s4_hselx,
  s4_hsize,
  s4_htrans,
  s4_hwdata,
  s4_hwrite,
  s5_haddr,
  s5_hburst,
  s5_hprot,
  s5_hrdata,
  s5_hready,
  s5_hresp,
  s5_hselx,
  s5_hsize,
  s5_htrans,
  s5_hwdata,
  s5_hwrite,
  s6_haddr,
  s6_hburst,
  s6_hprot,
  s6_hrdata,
  s6_hready,
  s6_hresp,
  s6_hselx,
  s6_hsize,
  s6_htrans,
  s6_hwdata,
  s6_hwrite,
  s7_haddr,
  s7_hburst,
  s7_hprot,
  s7_hrdata,
  s7_hready,
  s7_hresp,
  s7_hselx,
  s7_hsize,
  s7_htrans,
  s7_hwdata,
  s7_hwrite,
  s8_haddr,
  s8_hburst,
  s8_hprot,
  s8_hrdata,
  s8_hready,
  s8_hresp,
  s8_hselx,
  s8_hsize,
  s8_htrans,
  s8_hwdata,
  s8_hwrite,
  s9_haddr,
  s9_hburst,
  s9_hprot,
  s9_hrdata,
  s9_hready,
  s9_hresp,
  s9_hselx,
  s9_hsize,
  s9_htrans,
  s9_hwdata,
  s9_hwrite
);
input           hclk;           
input           hresetn;        
input   [31:0]  m0_haddr;       
input   [2 :0]  m0_hburst;      
input   [3 :0]  m0_hprot;       
input   [2 :0]  m0_hsize;       
input   [1 :0]  m0_htrans;      
input   [31:0]  m0_hwdata;      
input           m0_hwrite;      
input   [31:0]  m1_haddr;       
input   [2 :0]  m1_hburst;      
input   [3 :0]  m1_hprot;       
input   [2 :0]  m1_hsize;       
input   [1 :0]  m1_htrans;      
input   [31:0]  m1_hwdata;      
input           m1_hwrite;      
input   [31:0]  m2_haddr;       
input   [2 :0]  m2_hburst;      
input   [3 :0]  m2_hprot;       
input   [2 :0]  m2_hsize;       
input   [1 :0]  m2_htrans;      
input   [31:0]  m2_hwdata;      
input           m2_hwrite;      
input   [31:0]  m3_haddr;       
input   [2 :0]  m3_hburst;      
input   [3 :0]  m3_hprot;       
input   [2 :0]  m3_hsize;       
input   [1 :0]  m3_htrans;      
input   [31:0]  m3_hwdata;      
input           m3_hwrite;      
input   [31:0]  m4_haddr;       
input   [2 :0]  m4_hburst;      
input   [3 :0]  m4_hprot;       
input   [2 :0]  m4_hsize;       
input   [1 :0]  m4_htrans;      
input   [31:0]  m4_hwdata;      
input           m4_hwrite;      
input   [31:0]  m5_haddr;       
input   [2 :0]  m5_hburst;      
input   [3 :0]  m5_hprot;       
input   [2 :0]  m5_hsize;       
input   [1 :0]  m5_htrans;      
input   [31:0]  m5_hwdata;      
input           m5_hwrite;      
input   [31:0]  m6_haddr;       
input   [2 :0]  m6_hburst;      
input   [3 :0]  m6_hprot;       
input   [2 :0]  m6_hsize;       
input   [1 :0]  m6_htrans;      
input   [31:0]  m6_hwdata;      
input           m6_hwrite;      
input   [31:0]  s0_hrdata;      
input           s0_hready;      
input   [1 :0]  s0_hresp;       
input   [31:0]  s10_hrdata;     
input           s10_hready;     
input   [1 :0]  s10_hresp;      
input   [31:0]  s11_hrdata;     
input           s11_hready;     
input   [1 :0]  s11_hresp;      
input   [31:0]  s1_hrdata;      
input           s1_hready;      
input   [1 :0]  s1_hresp;       
input   [31:0]  s2_hrdata;      
input           s2_hready;      
input   [1 :0]  s2_hresp;       
input   [31:0]  s3_hrdata;      
input           s3_hready;      
input   [1 :0]  s3_hresp;       
input   [31:0]  s4_hrdata;      
input           s4_hready;      
input   [1 :0]  s4_hresp;       
input   [31:0]  s5_hrdata;      
input           s5_hready;      
input   [1 :0]  s5_hresp;       
input   [31:0]  s6_hrdata;      
input           s6_hready;      
input   [1 :0]  s6_hresp;       
input   [31:0]  s7_hrdata;      
input           s7_hready;      
input   [1 :0]  s7_hresp;       
input   [31:0]  s8_hrdata;      
input           s8_hready;      
input   [1 :0]  s8_hresp;       
input   [31:0]  s9_hrdata;      
input           s9_hready;      
input   [1 :0]  s9_hresp;       
output          m0_hgrant;      
output  [31:0]  m0_hrdata;      
output          m0_hready;      
output  [1 :0]  m0_hresp;       
output          m1_hgrant;      
output  [31:0]  m1_hrdata;      
output          m1_hready;      
output  [1 :0]  m1_hresp;       
output          m2_hgrant;      
output  [31:0]  m2_hrdata;      
output          m2_hready;      
output  [1 :0]  m2_hresp;       
output          m3_hgrant;      
output  [31:0]  m3_hrdata;      
output          m3_hready;      
output  [1 :0]  m3_hresp;       
output          m4_hgrant;      
output  [31:0]  m4_hrdata;      
output          m4_hready;      
output  [1 :0]  m4_hresp;       
output          m5_hgrant;      
output  [31:0]  m5_hrdata;      
output          m5_hready;      
output  [1 :0]  m5_hresp;       
output          m6_hgrant;      
output  [31:0]  m6_hrdata;      
output          m6_hready;      
output  [1 :0]  m6_hresp;       
output  [31:0]  s0_haddr;       
output  [2 :0]  s0_hburst;      
output  [3 :0]  s0_hprot;       
output          s0_hselx;       
output  [2 :0]  s0_hsize;       
output  [1 :0]  s0_htrans;      
output  [31:0]  s0_hwdata;      
output          s0_hwrite;      
output  [31:0]  s10_haddr;      
output  [2 :0]  s10_hburst;     
output  [3 :0]  s10_hprot;      
output          s10_hselx;      
output  [2 :0]  s10_hsize;      
output  [1 :0]  s10_htrans;     
output  [31:0]  s10_hwdata;     
output          s10_hwrite;     
output  [31:0]  s11_haddr;      
output  [2 :0]  s11_hburst;     
output  [3 :0]  s11_hprot;      
output          s11_hselx;      
output  [2 :0]  s11_hsize;      
output  [1 :0]  s11_htrans;     
output  [31:0]  s11_hwdata;     
output          s11_hwrite;     
output  [31:0]  s1_haddr;       
output  [2 :0]  s1_hburst;      
output  [3 :0]  s1_hprot;       
output          s1_hselx;       
output  [2 :0]  s1_hsize;       
output  [1 :0]  s1_htrans;      
output  [31:0]  s1_hwdata;      
output          s1_hwrite;      
output  [31:0]  s2_haddr;       
output  [2 :0]  s2_hburst;      
output  [3 :0]  s2_hprot;       
output          s2_hselx;       
output  [2 :0]  s2_hsize;       
output  [1 :0]  s2_htrans;      
output  [31:0]  s2_hwdata;      
output          s2_hwrite;      
output  [31:0]  s3_haddr;       
output  [2 :0]  s3_hburst;      
output  [3 :0]  s3_hprot;       
output          s3_hselx;       
output  [2 :0]  s3_hsize;       
output  [1 :0]  s3_htrans;      
output  [31:0]  s3_hwdata;      
output          s3_hwrite;      
output  [31:0]  s4_haddr;       
output  [2 :0]  s4_hburst;      
output  [3 :0]  s4_hprot;       
output          s4_hselx;       
output  [2 :0]  s4_hsize;       
output  [1 :0]  s4_htrans;      
output  [31:0]  s4_hwdata;      
output          s4_hwrite;      
output  [31:0]  s5_haddr;       
output  [2 :0]  s5_hburst;      
output  [3 :0]  s5_hprot;       
output          s5_hselx;       
output  [2 :0]  s5_hsize;       
output  [1 :0]  s5_htrans;      
output  [31:0]  s5_hwdata;      
output          s5_hwrite;      
output  [31:0]  s6_haddr;       
output  [2 :0]  s6_hburst;      
output  [3 :0]  s6_hprot;       
output          s6_hselx;       
output  [2 :0]  s6_hsize;       
output  [1 :0]  s6_htrans;      
output  [31:0]  s6_hwdata;      
output          s6_hwrite;      
output  [31:0]  s7_haddr;       
output  [2 :0]  s7_hburst;      
output  [3 :0]  s7_hprot;       
output          s7_hselx;       
output  [2 :0]  s7_hsize;       
output  [1 :0]  s7_htrans;      
output  [31:0]  s7_hwdata;      
output          s7_hwrite;      
output  [31:0]  s8_haddr;       
output  [2 :0]  s8_hburst;      
output  [3 :0]  s8_hprot;       
output          s8_hselx;       
output  [2 :0]  s8_hsize;       
output  [1 :0]  s8_htrans;      
output  [31:0]  s8_hwdata;      
output          s8_hwrite;      
output  [31:0]  s9_haddr;       
output  [2 :0]  s9_hburst;      
output  [3 :0]  s9_hprot;       
output          s9_hselx;       
output  [2 :0]  s9_hsize;       
output  [1 :0]  s9_htrans;      
output  [31:0]  s9_hwdata;      
output          s9_hwrite;      
wire            hclk;           
wire            hresetn;        
wire    [31:0]  m0_haddr;       
wire    [2 :0]  m0_hburst;      
wire            m0_hgrant;      
wire    [3 :0]  m0_hprot;       
wire    [31:0]  m0_hrdata;      
wire            m0_hready;      
wire    [1 :0]  m0_hresp;       
wire    [2 :0]  m0_hsize;       
wire    [1 :0]  m0_htrans;      
wire    [31:0]  m0_hwdata;      
wire            m0_hwrite;      
wire            m0_latch_cmd;   
wire            m0_nor_hready;  
wire            m0_s0_cmd_cur;  
wire            m0_s0_cmd_last; 
wire            m0_s0_data;     
wire            m0_s0_req;      
wire            m0_s10_cmd_cur; 
wire            m0_s10_cmd_last; 
wire            m0_s10_data;    
wire            m0_s10_req;     
wire            m0_s11_cmd_cur; 
wire            m0_s11_cmd_last; 
wire            m0_s11_data;    
wire            m0_s11_req;     
wire            m0_s1_cmd_cur;  
wire            m0_s1_cmd_last; 
wire            m0_s1_data;     
wire            m0_s1_req;      
wire            m0_s2_cmd_cur;  
wire            m0_s2_cmd_last; 
wire            m0_s2_data;     
wire            m0_s2_req;      
wire            m0_s3_cmd_cur;  
wire            m0_s3_cmd_last; 
wire            m0_s3_data;     
wire            m0_s3_req;      
wire            m0_s4_cmd_cur;  
wire            m0_s4_cmd_last; 
wire            m0_s4_data;     
wire            m0_s4_req;      
wire            m0_s5_cmd_cur;  
wire            m0_s5_cmd_last; 
wire            m0_s5_data;     
wire            m0_s5_req;      
wire            m0_s6_cmd_cur;  
wire            m0_s6_cmd_last; 
wire            m0_s6_data;     
wire            m0_s6_req;      
wire            m0_s7_cmd_cur;  
wire            m0_s7_cmd_last; 
wire            m0_s7_data;     
wire            m0_s7_req;      
wire            m0_s8_cmd_cur;  
wire            m0_s8_cmd_last; 
wire            m0_s8_data;     
wire            m0_s8_req;      
wire            m0_s9_cmd_cur;  
wire            m0_s9_cmd_last; 
wire            m0_s9_data;     
wire            m0_s9_req;      
wire    [31:0]  m1_haddr;       
wire    [2 :0]  m1_hburst;      
wire            m1_hgrant;      
wire    [3 :0]  m1_hprot;       
wire    [31:0]  m1_hrdata;      
wire            m1_hready;      
wire    [1 :0]  m1_hresp;       
wire    [2 :0]  m1_hsize;       
wire    [1 :0]  m1_htrans;      
wire    [31:0]  m1_hwdata;      
wire            m1_hwrite;      
wire            m1_latch_cmd;   
wire            m1_nor_hready;  
wire            m1_s0_cmd_cur;  
wire            m1_s0_cmd_last; 
wire            m1_s0_data;     
wire            m1_s0_req;      
wire            m1_s10_cmd_cur; 
wire            m1_s10_cmd_last; 
wire            m1_s10_data;    
wire            m1_s10_req;     
wire            m1_s11_cmd_cur; 
wire            m1_s11_cmd_last; 
wire            m1_s11_data;    
wire            m1_s11_req;     
wire            m1_s1_cmd_cur;  
wire            m1_s1_cmd_last; 
wire            m1_s1_data;     
wire            m1_s1_req;      
wire            m1_s2_cmd_cur;  
wire            m1_s2_cmd_last; 
wire            m1_s2_data;     
wire            m1_s2_req;      
wire            m1_s3_cmd_cur;  
wire            m1_s3_cmd_last; 
wire            m1_s3_data;     
wire            m1_s3_req;      
wire            m1_s4_cmd_cur;  
wire            m1_s4_cmd_last; 
wire            m1_s4_data;     
wire            m1_s4_req;      
wire            m1_s5_cmd_cur;  
wire            m1_s5_cmd_last; 
wire            m1_s5_data;     
wire            m1_s5_req;      
wire            m1_s6_cmd_cur;  
wire            m1_s6_cmd_last; 
wire            m1_s6_data;     
wire            m1_s6_req;      
wire            m1_s7_cmd_cur;  
wire            m1_s7_cmd_last; 
wire            m1_s7_data;     
wire            m1_s7_req;      
wire            m1_s8_cmd_cur;  
wire            m1_s8_cmd_last; 
wire            m1_s8_data;     
wire            m1_s8_req;      
wire            m1_s9_cmd_cur;  
wire            m1_s9_cmd_last; 
wire            m1_s9_data;     
wire            m1_s9_req;      
wire    [31:0]  m2_haddr;       
wire    [2 :0]  m2_hburst;      
wire            m2_hgrant;      
wire    [3 :0]  m2_hprot;       
wire    [31:0]  m2_hrdata;      
wire            m2_hready;      
wire    [1 :0]  m2_hresp;       
wire    [2 :0]  m2_hsize;       
wire    [1 :0]  m2_htrans;      
wire    [31:0]  m2_hwdata;      
wire            m2_hwrite;      
wire            m2_latch_cmd;   
wire            m2_nor_hready;  
wire            m2_s0_cmd_cur;  
wire            m2_s0_cmd_last; 
wire            m2_s0_data;     
wire            m2_s0_req;      
wire            m2_s10_cmd_cur; 
wire            m2_s10_cmd_last; 
wire            m2_s10_data;    
wire            m2_s10_req;     
wire            m2_s11_cmd_cur; 
wire            m2_s11_cmd_last; 
wire            m2_s11_data;    
wire            m2_s11_req;     
wire            m2_s1_cmd_cur;  
wire            m2_s1_cmd_last; 
wire            m2_s1_data;     
wire            m2_s1_req;      
wire            m2_s2_cmd_cur;  
wire            m2_s2_cmd_last; 
wire            m2_s2_data;     
wire            m2_s2_req;      
wire            m2_s3_cmd_cur;  
wire            m2_s3_cmd_last; 
wire            m2_s3_data;     
wire            m2_s3_req;      
wire            m2_s4_cmd_cur;  
wire            m2_s4_cmd_last; 
wire            m2_s4_data;     
wire            m2_s4_req;      
wire            m2_s5_cmd_cur;  
wire            m2_s5_cmd_last; 
wire            m2_s5_data;     
wire            m2_s5_req;      
wire            m2_s6_cmd_cur;  
wire            m2_s6_cmd_last; 
wire            m2_s6_data;     
wire            m2_s6_req;      
wire            m2_s7_cmd_cur;  
wire            m2_s7_cmd_last; 
wire            m2_s7_data;     
wire            m2_s7_req;      
wire            m2_s8_cmd_cur;  
wire            m2_s8_cmd_last; 
wire            m2_s8_data;     
wire            m2_s8_req;      
wire            m2_s9_cmd_cur;  
wire            m2_s9_cmd_last; 
wire            m2_s9_data;     
wire            m2_s9_req;      
wire    [31:0]  m3_haddr;       
wire    [2 :0]  m3_hburst;      
wire            m3_hgrant;      
wire    [3 :0]  m3_hprot;       
wire    [31:0]  m3_hrdata;      
wire            m3_hready;      
wire    [1 :0]  m3_hresp;       
wire    [2 :0]  m3_hsize;       
wire    [1 :0]  m3_htrans;      
wire    [31:0]  m3_hwdata;      
wire            m3_hwrite;      
wire            m3_latch_cmd;   
wire            m3_nor_hready;  
wire            m3_s0_cmd_cur;  
wire            m3_s0_cmd_last; 
wire            m3_s0_data;     
wire            m3_s0_req;      
wire            m3_s10_cmd_cur; 
wire            m3_s10_cmd_last; 
wire            m3_s10_data;    
wire            m3_s10_req;     
wire            m3_s11_cmd_cur; 
wire            m3_s11_cmd_last; 
wire            m3_s11_data;    
wire            m3_s11_req;     
wire            m3_s1_cmd_cur;  
wire            m3_s1_cmd_last; 
wire            m3_s1_data;     
wire            m3_s1_req;      
wire            m3_s2_cmd_cur;  
wire            m3_s2_cmd_last; 
wire            m3_s2_data;     
wire            m3_s2_req;      
wire            m3_s3_cmd_cur;  
wire            m3_s3_cmd_last; 
wire            m3_s3_data;     
wire            m3_s3_req;      
wire            m3_s4_cmd_cur;  
wire            m3_s4_cmd_last; 
wire            m3_s4_data;     
wire            m3_s4_req;      
wire            m3_s5_cmd_cur;  
wire            m3_s5_cmd_last; 
wire            m3_s5_data;     
wire            m3_s5_req;      
wire            m3_s6_cmd_cur;  
wire            m3_s6_cmd_last; 
wire            m3_s6_data;     
wire            m3_s6_req;      
wire            m3_s7_cmd_cur;  
wire            m3_s7_cmd_last; 
wire            m3_s7_data;     
wire            m3_s7_req;      
wire            m3_s8_cmd_cur;  
wire            m3_s8_cmd_last; 
wire            m3_s8_data;     
wire            m3_s8_req;      
wire            m3_s9_cmd_cur;  
wire            m3_s9_cmd_last; 
wire            m3_s9_data;     
wire            m3_s9_req;      
wire    [31:0]  m4_haddr;       
wire    [2 :0]  m4_hburst;      
wire            m4_hgrant;      
wire    [3 :0]  m4_hprot;       
wire    [31:0]  m4_hrdata;      
wire            m4_hready;      
wire    [1 :0]  m4_hresp;       
wire    [2 :0]  m4_hsize;       
wire    [1 :0]  m4_htrans;      
wire    [31:0]  m4_hwdata;      
wire            m4_hwrite;      
wire            m4_latch_cmd;   
wire            m4_nor_hready;  
wire            m4_s0_cmd_cur;  
wire            m4_s0_cmd_last; 
wire            m4_s0_data;     
wire            m4_s0_req;      
wire            m4_s10_cmd_cur; 
wire            m4_s10_cmd_last; 
wire            m4_s10_data;    
wire            m4_s10_req;     
wire            m4_s11_cmd_cur; 
wire            m4_s11_cmd_last; 
wire            m4_s11_data;    
wire            m4_s11_req;     
wire            m4_s1_cmd_cur;  
wire            m4_s1_cmd_last; 
wire            m4_s1_data;     
wire            m4_s1_req;      
wire            m4_s2_cmd_cur;  
wire            m4_s2_cmd_last; 
wire            m4_s2_data;     
wire            m4_s2_req;      
wire            m4_s3_cmd_cur;  
wire            m4_s3_cmd_last; 
wire            m4_s3_data;     
wire            m4_s3_req;      
wire            m4_s4_cmd_cur;  
wire            m4_s4_cmd_last; 
wire            m4_s4_data;     
wire            m4_s4_req;      
wire            m4_s5_cmd_cur;  
wire            m4_s5_cmd_last; 
wire            m4_s5_data;     
wire            m4_s5_req;      
wire            m4_s6_cmd_cur;  
wire            m4_s6_cmd_last; 
wire            m4_s6_data;     
wire            m4_s6_req;      
wire            m4_s7_cmd_cur;  
wire            m4_s7_cmd_last; 
wire            m4_s7_data;     
wire            m4_s7_req;      
wire            m4_s8_cmd_cur;  
wire            m4_s8_cmd_last; 
wire            m4_s8_data;     
wire            m4_s8_req;      
wire            m4_s9_cmd_cur;  
wire            m4_s9_cmd_last; 
wire            m4_s9_data;     
wire            m4_s9_req;      
wire    [31:0]  m5_haddr;       
wire    [2 :0]  m5_hburst;      
wire            m5_hgrant;      
wire    [3 :0]  m5_hprot;       
wire    [31:0]  m5_hrdata;      
wire            m5_hready;      
wire    [1 :0]  m5_hresp;       
wire    [2 :0]  m5_hsize;       
wire    [1 :0]  m5_htrans;      
wire    [31:0]  m5_hwdata;      
wire            m5_hwrite;      
wire            m5_latch_cmd;   
wire            m5_nor_hready;  
wire            m5_s0_cmd_cur;  
wire            m5_s0_cmd_last; 
wire            m5_s0_data;     
wire            m5_s0_req;      
wire            m5_s10_cmd_cur; 
wire            m5_s10_cmd_last; 
wire            m5_s10_data;    
wire            m5_s10_req;     
wire            m5_s11_cmd_cur; 
wire            m5_s11_cmd_last; 
wire            m5_s11_data;    
wire            m5_s11_req;     
wire            m5_s1_cmd_cur;  
wire            m5_s1_cmd_last; 
wire            m5_s1_data;     
wire            m5_s1_req;      
wire            m5_s2_cmd_cur;  
wire            m5_s2_cmd_last; 
wire            m5_s2_data;     
wire            m5_s2_req;      
wire            m5_s3_cmd_cur;  
wire            m5_s3_cmd_last; 
wire            m5_s3_data;     
wire            m5_s3_req;      
wire            m5_s4_cmd_cur;  
wire            m5_s4_cmd_last; 
wire            m5_s4_data;     
wire            m5_s4_req;      
wire            m5_s5_cmd_cur;  
wire            m5_s5_cmd_last; 
wire            m5_s5_data;     
wire            m5_s5_req;      
wire            m5_s6_cmd_cur;  
wire            m5_s6_cmd_last; 
wire            m5_s6_data;     
wire            m5_s6_req;      
wire            m5_s7_cmd_cur;  
wire            m5_s7_cmd_last; 
wire            m5_s7_data;     
wire            m5_s7_req;      
wire            m5_s8_cmd_cur;  
wire            m5_s8_cmd_last; 
wire            m5_s8_data;     
wire            m5_s8_req;      
wire            m5_s9_cmd_cur;  
wire            m5_s9_cmd_last; 
wire            m5_s9_data;     
wire            m5_s9_req;      
wire    [31:0]  m6_haddr;       
wire    [2 :0]  m6_hburst;      
wire            m6_hgrant;      
wire    [3 :0]  m6_hprot;       
wire    [31:0]  m6_hrdata;      
wire            m6_hready;      
wire    [1 :0]  m6_hresp;       
wire    [2 :0]  m6_hsize;       
wire    [1 :0]  m6_htrans;      
wire    [31:0]  m6_hwdata;      
wire            m6_hwrite;      
wire            m6_latch_cmd;   
wire            m6_nor_hready;  
wire            m6_s0_cmd_cur;  
wire            m6_s0_cmd_last; 
wire            m6_s0_data;     
wire            m6_s0_req;      
wire            m6_s10_cmd_cur; 
wire            m6_s10_cmd_last; 
wire            m6_s10_data;    
wire            m6_s10_req;     
wire            m6_s11_cmd_cur; 
wire            m6_s11_cmd_last; 
wire            m6_s11_data;    
wire            m6_s11_req;     
wire            m6_s1_cmd_cur;  
wire            m6_s1_cmd_last; 
wire            m6_s1_data;     
wire            m6_s1_req;      
wire            m6_s2_cmd_cur;  
wire            m6_s2_cmd_last; 
wire            m6_s2_data;     
wire            m6_s2_req;      
wire            m6_s3_cmd_cur;  
wire            m6_s3_cmd_last; 
wire            m6_s3_data;     
wire            m6_s3_req;      
wire            m6_s4_cmd_cur;  
wire            m6_s4_cmd_last; 
wire            m6_s4_data;     
wire            m6_s4_req;      
wire            m6_s5_cmd_cur;  
wire            m6_s5_cmd_last; 
wire            m6_s5_data;     
wire            m6_s5_req;      
wire            m6_s6_cmd_cur;  
wire            m6_s6_cmd_last; 
wire            m6_s6_data;     
wire            m6_s6_req;      
wire            m6_s7_cmd_cur;  
wire            m6_s7_cmd_last; 
wire            m6_s7_data;     
wire            m6_s7_req;      
wire            m6_s8_cmd_cur;  
wire            m6_s8_cmd_last; 
wire            m6_s8_data;     
wire            m6_s8_req;      
wire            m6_s9_cmd_cur;  
wire            m6_s9_cmd_last; 
wire            m6_s9_data;     
wire            m6_s9_req;      
wire    [31:0]  s0_haddr;       
wire    [2 :0]  s0_hburst;      
wire    [3 :0]  s0_hprot;       
wire    [31:0]  s0_hrdata;      
wire            s0_hready;      
wire    [1 :0]  s0_hresp;       
wire            s0_hselx;       
wire    [2 :0]  s0_hsize;       
wire    [1 :0]  s0_htrans;      
wire    [31:0]  s0_hwdata;      
wire            s0_hwrite;      
wire    [6 :0]  s0_req;         
wire    [31:0]  s10_haddr;      
wire    [2 :0]  s10_hburst;     
wire    [3 :0]  s10_hprot;      
wire    [31:0]  s10_hrdata;     
wire            s10_hready;     
wire    [1 :0]  s10_hresp;      
wire            s10_hselx;      
wire    [2 :0]  s10_hsize;      
wire    [1 :0]  s10_htrans;     
wire    [31:0]  s10_hwdata;     
wire            s10_hwrite;     
wire    [6 :0]  s10_req;        
wire    [31:0]  s11_haddr;      
wire    [2 :0]  s11_hburst;     
wire    [3 :0]  s11_hprot;      
wire    [31:0]  s11_hrdata;     
wire            s11_hready;     
wire    [1 :0]  s11_hresp;      
wire            s11_hselx;      
wire    [2 :0]  s11_hsize;      
wire    [1 :0]  s11_htrans;     
wire    [31:0]  s11_hwdata;     
wire            s11_hwrite;     
wire    [6 :0]  s11_req;        
wire    [31:0]  s1_haddr;       
wire    [2 :0]  s1_hburst;      
wire    [3 :0]  s1_hprot;       
wire    [31:0]  s1_hrdata;      
wire            s1_hready;      
wire    [1 :0]  s1_hresp;       
wire            s1_hselx;       
wire    [2 :0]  s1_hsize;       
wire    [1 :0]  s1_htrans;      
wire    [31:0]  s1_hwdata;      
wire            s1_hwrite;      
wire    [6 :0]  s1_req;         
wire    [31:0]  s2_haddr;       
wire    [2 :0]  s2_hburst;      
wire    [3 :0]  s2_hprot;       
wire    [31:0]  s2_hrdata;      
wire            s2_hready;      
wire    [1 :0]  s2_hresp;       
wire            s2_hselx;       
wire    [2 :0]  s2_hsize;       
wire    [1 :0]  s2_htrans;      
wire    [31:0]  s2_hwdata;      
wire            s2_hwrite;      
wire    [6 :0]  s2_req;         
wire    [31:0]  s3_haddr;       
wire    [2 :0]  s3_hburst;      
wire    [3 :0]  s3_hprot;       
wire    [31:0]  s3_hrdata;      
wire            s3_hready;      
wire    [1 :0]  s3_hresp;       
wire            s3_hselx;       
wire    [2 :0]  s3_hsize;       
wire    [1 :0]  s3_htrans;      
wire    [31:0]  s3_hwdata;      
wire            s3_hwrite;      
wire    [6 :0]  s3_req;         
wire    [31:0]  s4_haddr;       
wire    [2 :0]  s4_hburst;      
wire    [3 :0]  s4_hprot;       
wire    [31:0]  s4_hrdata;      
wire            s4_hready;      
wire    [1 :0]  s4_hresp;       
wire            s4_hselx;       
wire    [2 :0]  s4_hsize;       
wire    [1 :0]  s4_htrans;      
wire    [31:0]  s4_hwdata;      
wire            s4_hwrite;      
wire    [6 :0]  s4_req;         
wire    [31:0]  s5_haddr;       
wire    [2 :0]  s5_hburst;      
wire    [3 :0]  s5_hprot;       
wire    [31:0]  s5_hrdata;      
wire            s5_hready;      
wire    [1 :0]  s5_hresp;       
wire            s5_hselx;       
wire    [2 :0]  s5_hsize;       
wire    [1 :0]  s5_htrans;      
wire    [31:0]  s5_hwdata;      
wire            s5_hwrite;      
wire    [6 :0]  s5_req;         
wire    [31:0]  s6_haddr;       
wire    [2 :0]  s6_hburst;      
wire    [3 :0]  s6_hprot;       
wire    [31:0]  s6_hrdata;      
wire            s6_hready;      
wire    [1 :0]  s6_hresp;       
wire            s6_hselx;       
wire    [2 :0]  s6_hsize;       
wire    [1 :0]  s6_htrans;      
wire    [31:0]  s6_hwdata;      
wire            s6_hwrite;      
wire    [6 :0]  s6_req;         
wire    [31:0]  s7_haddr;       
wire    [2 :0]  s7_hburst;      
wire    [3 :0]  s7_hprot;       
wire    [31:0]  s7_hrdata;      
wire            s7_hready;      
wire    [1 :0]  s7_hresp;       
wire            s7_hselx;       
wire    [2 :0]  s7_hsize;       
wire    [1 :0]  s7_htrans;      
wire    [31:0]  s7_hwdata;      
wire            s7_hwrite;      
wire    [6 :0]  s7_req;         
wire    [31:0]  s8_haddr;       
wire    [2 :0]  s8_hburst;      
wire    [3 :0]  s8_hprot;       
wire    [31:0]  s8_hrdata;      
wire            s8_hready;      
wire    [1 :0]  s8_hresp;       
wire            s8_hselx;       
wire    [2 :0]  s8_hsize;       
wire    [1 :0]  s8_htrans;      
wire    [31:0]  s8_hwdata;      
wire            s8_hwrite;      
wire    [6 :0]  s8_req;         
wire    [31:0]  s9_haddr;       
wire    [2 :0]  s9_hburst;      
wire    [3 :0]  s9_hprot;       
wire    [31:0]  s9_hrdata;      
wire            s9_hready;      
wire    [1 :0]  s9_hresp;       
wire            s9_hselx;       
wire    [2 :0]  s9_hsize;       
wire    [1 :0]  s9_htrans;      
wire    [31:0]  s9_hwdata;      
wire            s9_hwrite;      
wire    [6 :0]  s9_req;         
ahb_matrix_7_12_dec  x_matrix_dec (
  .hclk            (hclk           ),
  .hresetn         (hresetn        ),
  .m0_haddr        (m0_haddr       ),
  .m0_hburst       (m0_hburst      ),
  .m0_hgrant       (m0_hgrant      ),
  .m0_hprot        (m0_hprot       ),
  .m0_hrdata       (m0_hrdata      ),
  .m0_hready       (m0_hready      ),
  .m0_hresp        (m0_hresp       ),
  .m0_hsize        (m0_hsize       ),
  .m0_htrans       (m0_htrans      ),
  .m0_hwdata       (m0_hwdata      ),
  .m0_hwrite       (m0_hwrite      ),
  .m0_latch_cmd    (m0_latch_cmd   ),
  .m0_nor_hready   (m0_nor_hready  ),
  .m0_s0_cmd_cur   (m0_s0_cmd_cur  ),
  .m0_s0_cmd_last  (m0_s0_cmd_last ),
  .m0_s0_data      (m0_s0_data     ),
  .m0_s0_req       (m0_s0_req      ),
  .m0_s10_cmd_cur  (m0_s10_cmd_cur ),
  .m0_s10_cmd_last (m0_s10_cmd_last),
  .m0_s10_data     (m0_s10_data    ),
  .m0_s10_req      (m0_s10_req     ),
  .m0_s11_cmd_cur  (m0_s11_cmd_cur ),
  .m0_s11_cmd_last (m0_s11_cmd_last),
  .m0_s11_data     (m0_s11_data    ),
  .m0_s11_req      (m0_s11_req     ),
  .m0_s1_cmd_cur   (m0_s1_cmd_cur  ),
  .m0_s1_cmd_last  (m0_s1_cmd_last ),
  .m0_s1_data      (m0_s1_data     ),
  .m0_s1_req       (m0_s1_req      ),
  .m0_s2_cmd_cur   (m0_s2_cmd_cur  ),
  .m0_s2_cmd_last  (m0_s2_cmd_last ),
  .m0_s2_data      (m0_s2_data     ),
  .m0_s2_req       (m0_s2_req      ),
  .m0_s3_cmd_cur   (m0_s3_cmd_cur  ),
  .m0_s3_cmd_last  (m0_s3_cmd_last ),
  .m0_s3_data      (m0_s3_data     ),
  .m0_s3_req       (m0_s3_req      ),
  .m0_s4_cmd_cur   (m0_s4_cmd_cur  ),
  .m0_s4_cmd_last  (m0_s4_cmd_last ),
  .m0_s4_data      (m0_s4_data     ),
  .m0_s4_req       (m0_s4_req      ),
  .m0_s5_cmd_cur   (m0_s5_cmd_cur  ),
  .m0_s5_cmd_last  (m0_s5_cmd_last ),
  .m0_s5_data      (m0_s5_data     ),
  .m0_s5_req       (m0_s5_req      ),
  .m0_s6_cmd_cur   (m0_s6_cmd_cur  ),
  .m0_s6_cmd_last  (m0_s6_cmd_last ),
  .m0_s6_data      (m0_s6_data     ),
  .m0_s6_req       (m0_s6_req      ),
  .m0_s7_cmd_cur   (m0_s7_cmd_cur  ),
  .m0_s7_cmd_last  (m0_s7_cmd_last ),
  .m0_s7_data      (m0_s7_data     ),
  .m0_s7_req       (m0_s7_req      ),
  .m0_s8_cmd_cur   (m0_s8_cmd_cur  ),
  .m0_s8_cmd_last  (m0_s8_cmd_last ),
  .m0_s8_data      (m0_s8_data     ),
  .m0_s8_req       (m0_s8_req      ),
  .m0_s9_cmd_cur   (m0_s9_cmd_cur  ),
  .m0_s9_cmd_last  (m0_s9_cmd_last ),
  .m0_s9_data      (m0_s9_data     ),
  .m0_s9_req       (m0_s9_req      ),
  .m1_haddr        (m1_haddr       ),
  .m1_hburst       (m1_hburst      ),
  .m1_hgrant       (m1_hgrant      ),
  .m1_hprot        (m1_hprot       ),
  .m1_hrdata       (m1_hrdata      ),
  .m1_hready       (m1_hready      ),
  .m1_hresp        (m1_hresp       ),
  .m1_hsize        (m1_hsize       ),
  .m1_htrans       (m1_htrans      ),
  .m1_hwdata       (m1_hwdata      ),
  .m1_hwrite       (m1_hwrite      ),
  .m1_latch_cmd    (m1_latch_cmd   ),
  .m1_nor_hready   (m1_nor_hready  ),
  .m1_s0_cmd_cur   (m1_s0_cmd_cur  ),
  .m1_s0_cmd_last  (m1_s0_cmd_last ),
  .m1_s0_data      (m1_s0_data     ),
  .m1_s0_req       (m1_s0_req      ),
  .m1_s10_cmd_cur  (m1_s10_cmd_cur ),
  .m1_s10_cmd_last (m1_s10_cmd_last),
  .m1_s10_data     (m1_s10_data    ),
  .m1_s10_req      (m1_s10_req     ),
  .m1_s11_cmd_cur  (m1_s11_cmd_cur ),
  .m1_s11_cmd_last (m1_s11_cmd_last),
  .m1_s11_data     (m1_s11_data    ),
  .m1_s11_req      (m1_s11_req     ),
  .m1_s1_cmd_cur   (m1_s1_cmd_cur  ),
  .m1_s1_cmd_last  (m1_s1_cmd_last ),
  .m1_s1_data      (m1_s1_data     ),
  .m1_s1_req       (m1_s1_req      ),
  .m1_s2_cmd_cur   (m1_s2_cmd_cur  ),
  .m1_s2_cmd_last  (m1_s2_cmd_last ),
  .m1_s2_data      (m1_s2_data     ),
  .m1_s2_req       (m1_s2_req      ),
  .m1_s3_cmd_cur   (m1_s3_cmd_cur  ),
  .m1_s3_cmd_last  (m1_s3_cmd_last ),
  .m1_s3_data      (m1_s3_data     ),
  .m1_s3_req       (m1_s3_req      ),
  .m1_s4_cmd_cur   (m1_s4_cmd_cur  ),
  .m1_s4_cmd_last  (m1_s4_cmd_last ),
  .m1_s4_data      (m1_s4_data     ),
  .m1_s4_req       (m1_s4_req      ),
  .m1_s5_cmd_cur   (m1_s5_cmd_cur  ),
  .m1_s5_cmd_last  (m1_s5_cmd_last ),
  .m1_s5_data      (m1_s5_data     ),
  .m1_s5_req       (m1_s5_req      ),
  .m1_s6_cmd_cur   (m1_s6_cmd_cur  ),
  .m1_s6_cmd_last  (m1_s6_cmd_last ),
  .m1_s6_data      (m1_s6_data     ),
  .m1_s6_req       (m1_s6_req      ),
  .m1_s7_cmd_cur   (m1_s7_cmd_cur  ),
  .m1_s7_cmd_last  (m1_s7_cmd_last ),
  .m1_s7_data      (m1_s7_data     ),
  .m1_s7_req       (m1_s7_req      ),
  .m1_s8_cmd_cur   (m1_s8_cmd_cur  ),
  .m1_s8_cmd_last  (m1_s8_cmd_last ),
  .m1_s8_data      (m1_s8_data     ),
  .m1_s8_req       (m1_s8_req      ),
  .m1_s9_cmd_cur   (m1_s9_cmd_cur  ),
  .m1_s9_cmd_last  (m1_s9_cmd_last ),
  .m1_s9_data      (m1_s9_data     ),
  .m1_s9_req       (m1_s9_req      ),
  .m2_haddr        (m2_haddr       ),
  .m2_hburst       (m2_hburst      ),
  .m2_hgrant       (m2_hgrant      ),
  .m2_hprot        (m2_hprot       ),
  .m2_hrdata       (m2_hrdata      ),
  .m2_hready       (m2_hready      ),
  .m2_hresp        (m2_hresp       ),
  .m2_hsize        (m2_hsize       ),
  .m2_htrans       (m2_htrans      ),
  .m2_hwdata       (m2_hwdata      ),
  .m2_hwrite       (m2_hwrite      ),
  .m2_latch_cmd    (m2_latch_cmd   ),
  .m2_nor_hready   (m2_nor_hready  ),
  .m2_s0_cmd_cur   (m2_s0_cmd_cur  ),
  .m2_s0_cmd_last  (m2_s0_cmd_last ),
  .m2_s0_data      (m2_s0_data     ),
  .m2_s0_req       (m2_s0_req      ),
  .m2_s10_cmd_cur  (m2_s10_cmd_cur ),
  .m2_s10_cmd_last (m2_s10_cmd_last),
  .m2_s10_data     (m2_s10_data    ),
  .m2_s10_req      (m2_s10_req     ),
  .m2_s11_cmd_cur  (m2_s11_cmd_cur ),
  .m2_s11_cmd_last (m2_s11_cmd_last),
  .m2_s11_data     (m2_s11_data    ),
  .m2_s11_req      (m2_s11_req     ),
  .m2_s1_cmd_cur   (m2_s1_cmd_cur  ),
  .m2_s1_cmd_last  (m2_s1_cmd_last ),
  .m2_s1_data      (m2_s1_data     ),
  .m2_s1_req       (m2_s1_req      ),
  .m2_s2_cmd_cur   (m2_s2_cmd_cur  ),
  .m2_s2_cmd_last  (m2_s2_cmd_last ),
  .m2_s2_data      (m2_s2_data     ),
  .m2_s2_req       (m2_s2_req      ),
  .m2_s3_cmd_cur   (m2_s3_cmd_cur  ),
  .m2_s3_cmd_last  (m2_s3_cmd_last ),
  .m2_s3_data      (m2_s3_data     ),
  .m2_s3_req       (m2_s3_req      ),
  .m2_s4_cmd_cur   (m2_s4_cmd_cur  ),
  .m2_s4_cmd_last  (m2_s4_cmd_last ),
  .m2_s4_data      (m2_s4_data     ),
  .m2_s4_req       (m2_s4_req      ),
  .m2_s5_cmd_cur   (m2_s5_cmd_cur  ),
  .m2_s5_cmd_last  (m2_s5_cmd_last ),
  .m2_s5_data      (m2_s5_data     ),
  .m2_s5_req       (m2_s5_req      ),
  .m2_s6_cmd_cur   (m2_s6_cmd_cur  ),
  .m2_s6_cmd_last  (m2_s6_cmd_last ),
  .m2_s6_data      (m2_s6_data     ),
  .m2_s6_req       (m2_s6_req      ),
  .m2_s7_cmd_cur   (m2_s7_cmd_cur  ),
  .m2_s7_cmd_last  (m2_s7_cmd_last ),
  .m2_s7_data      (m2_s7_data     ),
  .m2_s7_req       (m2_s7_req      ),
  .m2_s8_cmd_cur   (m2_s8_cmd_cur  ),
  .m2_s8_cmd_last  (m2_s8_cmd_last ),
  .m2_s8_data      (m2_s8_data     ),
  .m2_s8_req       (m2_s8_req      ),
  .m2_s9_cmd_cur   (m2_s9_cmd_cur  ),
  .m2_s9_cmd_last  (m2_s9_cmd_last ),
  .m2_s9_data      (m2_s9_data     ),
  .m2_s9_req       (m2_s9_req      ),
  .m3_haddr        (m3_haddr       ),
  .m3_hburst       (m3_hburst      ),
  .m3_hgrant       (m3_hgrant      ),
  .m3_hprot        (m3_hprot       ),
  .m3_hrdata       (m3_hrdata      ),
  .m3_hready       (m3_hready      ),
  .m3_hresp        (m3_hresp       ),
  .m3_hsize        (m3_hsize       ),
  .m3_htrans       (m3_htrans      ),
  .m3_hwdata       (m3_hwdata      ),
  .m3_hwrite       (m3_hwrite      ),
  .m3_latch_cmd    (m3_latch_cmd   ),
  .m3_nor_hready   (m3_nor_hready  ),
  .m3_s0_cmd_cur   (m3_s0_cmd_cur  ),
  .m3_s0_cmd_last  (m3_s0_cmd_last ),
  .m3_s0_data      (m3_s0_data     ),
  .m3_s0_req       (m3_s0_req      ),
  .m3_s10_cmd_cur  (m3_s10_cmd_cur ),
  .m3_s10_cmd_last (m3_s10_cmd_last),
  .m3_s10_data     (m3_s10_data    ),
  .m3_s10_req      (m3_s10_req     ),
  .m3_s11_cmd_cur  (m3_s11_cmd_cur ),
  .m3_s11_cmd_last (m3_s11_cmd_last),
  .m3_s11_data     (m3_s11_data    ),
  .m3_s11_req      (m3_s11_req     ),
  .m3_s1_cmd_cur   (m3_s1_cmd_cur  ),
  .m3_s1_cmd_last  (m3_s1_cmd_last ),
  .m3_s1_data      (m3_s1_data     ),
  .m3_s1_req       (m3_s1_req      ),
  .m3_s2_cmd_cur   (m3_s2_cmd_cur  ),
  .m3_s2_cmd_last  (m3_s2_cmd_last ),
  .m3_s2_data      (m3_s2_data     ),
  .m3_s2_req       (m3_s2_req      ),
  .m3_s3_cmd_cur   (m3_s3_cmd_cur  ),
  .m3_s3_cmd_last  (m3_s3_cmd_last ),
  .m3_s3_data      (m3_s3_data     ),
  .m3_s3_req       (m3_s3_req      ),
  .m3_s4_cmd_cur   (m3_s4_cmd_cur  ),
  .m3_s4_cmd_last  (m3_s4_cmd_last ),
  .m3_s4_data      (m3_s4_data     ),
  .m3_s4_req       (m3_s4_req      ),
  .m3_s5_cmd_cur   (m3_s5_cmd_cur  ),
  .m3_s5_cmd_last  (m3_s5_cmd_last ),
  .m3_s5_data      (m3_s5_data     ),
  .m3_s5_req       (m3_s5_req      ),
  .m3_s6_cmd_cur   (m3_s6_cmd_cur  ),
  .m3_s6_cmd_last  (m3_s6_cmd_last ),
  .m3_s6_data      (m3_s6_data     ),
  .m3_s6_req       (m3_s6_req      ),
  .m3_s7_cmd_cur   (m3_s7_cmd_cur  ),
  .m3_s7_cmd_last  (m3_s7_cmd_last ),
  .m3_s7_data      (m3_s7_data     ),
  .m3_s7_req       (m3_s7_req      ),
  .m3_s8_cmd_cur   (m3_s8_cmd_cur  ),
  .m3_s8_cmd_last  (m3_s8_cmd_last ),
  .m3_s8_data      (m3_s8_data     ),
  .m3_s8_req       (m3_s8_req      ),
  .m3_s9_cmd_cur   (m3_s9_cmd_cur  ),
  .m3_s9_cmd_last  (m3_s9_cmd_last ),
  .m3_s9_data      (m3_s9_data     ),
  .m3_s9_req       (m3_s9_req      ),
  .m4_haddr        (m4_haddr       ),
  .m4_hburst       (m4_hburst      ),
  .m4_hgrant       (m4_hgrant      ),
  .m4_hprot        (m4_hprot       ),
  .m4_hrdata       (m4_hrdata      ),
  .m4_hready       (m4_hready      ),
  .m4_hresp        (m4_hresp       ),
  .m4_hsize        (m4_hsize       ),
  .m4_htrans       (m4_htrans      ),
  .m4_hwdata       (m4_hwdata      ),
  .m4_hwrite       (m4_hwrite      ),
  .m4_latch_cmd    (m4_latch_cmd   ),
  .m4_nor_hready   (m4_nor_hready  ),
  .m4_s0_cmd_cur   (m4_s0_cmd_cur  ),
  .m4_s0_cmd_last  (m4_s0_cmd_last ),
  .m4_s0_data      (m4_s0_data     ),
  .m4_s0_req       (m4_s0_req      ),
  .m4_s10_cmd_cur  (m4_s10_cmd_cur ),
  .m4_s10_cmd_last (m4_s10_cmd_last),
  .m4_s10_data     (m4_s10_data    ),
  .m4_s10_req      (m4_s10_req     ),
  .m4_s11_cmd_cur  (m4_s11_cmd_cur ),
  .m4_s11_cmd_last (m4_s11_cmd_last),
  .m4_s11_data     (m4_s11_data    ),
  .m4_s11_req      (m4_s11_req     ),
  .m4_s1_cmd_cur   (m4_s1_cmd_cur  ),
  .m4_s1_cmd_last  (m4_s1_cmd_last ),
  .m4_s1_data      (m4_s1_data     ),
  .m4_s1_req       (m4_s1_req      ),
  .m4_s2_cmd_cur   (m4_s2_cmd_cur  ),
  .m4_s2_cmd_last  (m4_s2_cmd_last ),
  .m4_s2_data      (m4_s2_data     ),
  .m4_s2_req       (m4_s2_req      ),
  .m4_s3_cmd_cur   (m4_s3_cmd_cur  ),
  .m4_s3_cmd_last  (m4_s3_cmd_last ),
  .m4_s3_data      (m4_s3_data     ),
  .m4_s3_req       (m4_s3_req      ),
  .m4_s4_cmd_cur   (m4_s4_cmd_cur  ),
  .m4_s4_cmd_last  (m4_s4_cmd_last ),
  .m4_s4_data      (m4_s4_data     ),
  .m4_s4_req       (m4_s4_req      ),
  .m4_s5_cmd_cur   (m4_s5_cmd_cur  ),
  .m4_s5_cmd_last  (m4_s5_cmd_last ),
  .m4_s5_data      (m4_s5_data     ),
  .m4_s5_req       (m4_s5_req      ),
  .m4_s6_cmd_cur   (m4_s6_cmd_cur  ),
  .m4_s6_cmd_last  (m4_s6_cmd_last ),
  .m4_s6_data      (m4_s6_data     ),
  .m4_s6_req       (m4_s6_req      ),
  .m4_s7_cmd_cur   (m4_s7_cmd_cur  ),
  .m4_s7_cmd_last  (m4_s7_cmd_last ),
  .m4_s7_data      (m4_s7_data     ),
  .m4_s7_req       (m4_s7_req      ),
  .m4_s8_cmd_cur   (m4_s8_cmd_cur  ),
  .m4_s8_cmd_last  (m4_s8_cmd_last ),
  .m4_s8_data      (m4_s8_data     ),
  .m4_s8_req       (m4_s8_req      ),
  .m4_s9_cmd_cur   (m4_s9_cmd_cur  ),
  .m4_s9_cmd_last  (m4_s9_cmd_last ),
  .m4_s9_data      (m4_s9_data     ),
  .m4_s9_req       (m4_s9_req      ),
  .m5_haddr        (m5_haddr       ),
  .m5_hburst       (m5_hburst      ),
  .m5_hgrant       (m5_hgrant      ),
  .m5_hprot        (m5_hprot       ),
  .m5_hrdata       (m5_hrdata      ),
  .m5_hready       (m5_hready      ),
  .m5_hresp        (m5_hresp       ),
  .m5_hsize        (m5_hsize       ),
  .m5_htrans       (m5_htrans      ),
  .m5_hwdata       (m5_hwdata      ),
  .m5_hwrite       (m5_hwrite      ),
  .m5_latch_cmd    (m5_latch_cmd   ),
  .m5_nor_hready   (m5_nor_hready  ),
  .m5_s0_cmd_cur   (m5_s0_cmd_cur  ),
  .m5_s0_cmd_last  (m5_s0_cmd_last ),
  .m5_s0_data      (m5_s0_data     ),
  .m5_s0_req       (m5_s0_req      ),
  .m5_s10_cmd_cur  (m5_s10_cmd_cur ),
  .m5_s10_cmd_last (m5_s10_cmd_last),
  .m5_s10_data     (m5_s10_data    ),
  .m5_s10_req      (m5_s10_req     ),
  .m5_s11_cmd_cur  (m5_s11_cmd_cur ),
  .m5_s11_cmd_last (m5_s11_cmd_last),
  .m5_s11_data     (m5_s11_data    ),
  .m5_s11_req      (m5_s11_req     ),
  .m5_s1_cmd_cur   (m5_s1_cmd_cur  ),
  .m5_s1_cmd_last  (m5_s1_cmd_last ),
  .m5_s1_data      (m5_s1_data     ),
  .m5_s1_req       (m5_s1_req      ),
  .m5_s2_cmd_cur   (m5_s2_cmd_cur  ),
  .m5_s2_cmd_last  (m5_s2_cmd_last ),
  .m5_s2_data      (m5_s2_data     ),
  .m5_s2_req       (m5_s2_req      ),
  .m5_s3_cmd_cur   (m5_s3_cmd_cur  ),
  .m5_s3_cmd_last  (m5_s3_cmd_last ),
  .m5_s3_data      (m5_s3_data     ),
  .m5_s3_req       (m5_s3_req      ),
  .m5_s4_cmd_cur   (m5_s4_cmd_cur  ),
  .m5_s4_cmd_last  (m5_s4_cmd_last ),
  .m5_s4_data      (m5_s4_data     ),
  .m5_s4_req       (m5_s4_req      ),
  .m5_s5_cmd_cur   (m5_s5_cmd_cur  ),
  .m5_s5_cmd_last  (m5_s5_cmd_last ),
  .m5_s5_data      (m5_s5_data     ),
  .m5_s5_req       (m5_s5_req      ),
  .m5_s6_cmd_cur   (m5_s6_cmd_cur  ),
  .m5_s6_cmd_last  (m5_s6_cmd_last ),
  .m5_s6_data      (m5_s6_data     ),
  .m5_s6_req       (m5_s6_req      ),
  .m5_s7_cmd_cur   (m5_s7_cmd_cur  ),
  .m5_s7_cmd_last  (m5_s7_cmd_last ),
  .m5_s7_data      (m5_s7_data     ),
  .m5_s7_req       (m5_s7_req      ),
  .m5_s8_cmd_cur   (m5_s8_cmd_cur  ),
  .m5_s8_cmd_last  (m5_s8_cmd_last ),
  .m5_s8_data      (m5_s8_data     ),
  .m5_s8_req       (m5_s8_req      ),
  .m5_s9_cmd_cur   (m5_s9_cmd_cur  ),
  .m5_s9_cmd_last  (m5_s9_cmd_last ),
  .m5_s9_data      (m5_s9_data     ),
  .m5_s9_req       (m5_s9_req      ),
  .m6_haddr        (m6_haddr       ),
  .m6_hburst       (m6_hburst      ),
  .m6_hgrant       (m6_hgrant      ),
  .m6_hprot        (m6_hprot       ),
  .m6_hrdata       (m6_hrdata      ),
  .m6_hready       (m6_hready      ),
  .m6_hresp        (m6_hresp       ),
  .m6_hsize        (m6_hsize       ),
  .m6_htrans       (m6_htrans      ),
  .m6_hwdata       (m6_hwdata      ),
  .m6_hwrite       (m6_hwrite      ),
  .m6_latch_cmd    (m6_latch_cmd   ),
  .m6_nor_hready   (m6_nor_hready  ),
  .m6_s0_cmd_cur   (m6_s0_cmd_cur  ),
  .m6_s0_cmd_last  (m6_s0_cmd_last ),
  .m6_s0_data      (m6_s0_data     ),
  .m6_s0_req       (m6_s0_req      ),
  .m6_s10_cmd_cur  (m6_s10_cmd_cur ),
  .m6_s10_cmd_last (m6_s10_cmd_last),
  .m6_s10_data     (m6_s10_data    ),
  .m6_s10_req      (m6_s10_req     ),
  .m6_s11_cmd_cur  (m6_s11_cmd_cur ),
  .m6_s11_cmd_last (m6_s11_cmd_last),
  .m6_s11_data     (m6_s11_data    ),
  .m6_s11_req      (m6_s11_req     ),
  .m6_s1_cmd_cur   (m6_s1_cmd_cur  ),
  .m6_s1_cmd_last  (m6_s1_cmd_last ),
  .m6_s1_data      (m6_s1_data     ),
  .m6_s1_req       (m6_s1_req      ),
  .m6_s2_cmd_cur   (m6_s2_cmd_cur  ),
  .m6_s2_cmd_last  (m6_s2_cmd_last ),
  .m6_s2_data      (m6_s2_data     ),
  .m6_s2_req       (m6_s2_req      ),
  .m6_s3_cmd_cur   (m6_s3_cmd_cur  ),
  .m6_s3_cmd_last  (m6_s3_cmd_last ),
  .m6_s3_data      (m6_s3_data     ),
  .m6_s3_req       (m6_s3_req      ),
  .m6_s4_cmd_cur   (m6_s4_cmd_cur  ),
  .m6_s4_cmd_last  (m6_s4_cmd_last ),
  .m6_s4_data      (m6_s4_data     ),
  .m6_s4_req       (m6_s4_req      ),
  .m6_s5_cmd_cur   (m6_s5_cmd_cur  ),
  .m6_s5_cmd_last  (m6_s5_cmd_last ),
  .m6_s5_data      (m6_s5_data     ),
  .m6_s5_req       (m6_s5_req      ),
  .m6_s6_cmd_cur   (m6_s6_cmd_cur  ),
  .m6_s6_cmd_last  (m6_s6_cmd_last ),
  .m6_s6_data      (m6_s6_data     ),
  .m6_s6_req       (m6_s6_req      ),
  .m6_s7_cmd_cur   (m6_s7_cmd_cur  ),
  .m6_s7_cmd_last  (m6_s7_cmd_last ),
  .m6_s7_data      (m6_s7_data     ),
  .m6_s7_req       (m6_s7_req      ),
  .m6_s8_cmd_cur   (m6_s8_cmd_cur  ),
  .m6_s8_cmd_last  (m6_s8_cmd_last ),
  .m6_s8_data      (m6_s8_data     ),
  .m6_s8_req       (m6_s8_req      ),
  .m6_s9_cmd_cur   (m6_s9_cmd_cur  ),
  .m6_s9_cmd_last  (m6_s9_cmd_last ),
  .m6_s9_data      (m6_s9_data     ),
  .m6_s9_req       (m6_s9_req      ),
  .s0_haddr        (s0_haddr       ),
  .s0_hburst       (s0_hburst      ),
  .s0_hprot        (s0_hprot       ),
  .s0_hrdata       (s0_hrdata      ),
  .s0_hresp        (s0_hresp       ),
  .s0_hselx        (s0_hselx       ),
  .s0_hsize        (s0_hsize       ),
  .s0_htrans       (s0_htrans      ),
  .s0_hwdata       (s0_hwdata      ),
  .s0_hwrite       (s0_hwrite      ),
  .s0_req          (s0_req         ),
  .s10_haddr       (s10_haddr      ),
  .s10_hburst      (s10_hburst     ),
  .s10_hprot       (s10_hprot      ),
  .s10_hrdata      (s10_hrdata     ),
  .s10_hresp       (s10_hresp      ),
  .s10_hselx       (s10_hselx      ),
  .s10_hsize       (s10_hsize      ),
  .s10_htrans      (s10_htrans     ),
  .s10_hwdata      (s10_hwdata     ),
  .s10_hwrite      (s10_hwrite     ),
  .s10_req         (s10_req        ),
  .s11_haddr       (s11_haddr      ),
  .s11_hburst      (s11_hburst     ),
  .s11_hprot       (s11_hprot      ),
  .s11_hrdata      (s11_hrdata     ),
  .s11_hresp       (s11_hresp      ),
  .s11_hselx       (s11_hselx      ),
  .s11_hsize       (s11_hsize      ),
  .s11_htrans      (s11_htrans     ),
  .s11_hwdata      (s11_hwdata     ),
  .s11_hwrite      (s11_hwrite     ),
  .s11_req         (s11_req        ),
  .s1_haddr        (s1_haddr       ),
  .s1_hburst       (s1_hburst      ),
  .s1_hprot        (s1_hprot       ),
  .s1_hrdata       (s1_hrdata      ),
  .s1_hresp        (s1_hresp       ),
  .s1_hselx        (s1_hselx       ),
  .s1_hsize        (s1_hsize       ),
  .s1_htrans       (s1_htrans      ),
  .s1_hwdata       (s1_hwdata      ),
  .s1_hwrite       (s1_hwrite      ),
  .s1_req          (s1_req         ),
  .s2_haddr        (s2_haddr       ),
  .s2_hburst       (s2_hburst      ),
  .s2_hprot        (s2_hprot       ),
  .s2_hrdata       (s2_hrdata      ),
  .s2_hresp        (s2_hresp       ),
  .s2_hselx        (s2_hselx       ),
  .s2_hsize        (s2_hsize       ),
  .s2_htrans       (s2_htrans      ),
  .s2_hwdata       (s2_hwdata      ),
  .s2_hwrite       (s2_hwrite      ),
  .s2_req          (s2_req         ),
  .s3_haddr        (s3_haddr       ),
  .s3_hburst       (s3_hburst      ),
  .s3_hprot        (s3_hprot       ),
  .s3_hrdata       (s3_hrdata      ),
  .s3_hresp        (s3_hresp       ),
  .s3_hselx        (s3_hselx       ),
  .s3_hsize        (s3_hsize       ),
  .s3_htrans       (s3_htrans      ),
  .s3_hwdata       (s3_hwdata      ),
  .s3_hwrite       (s3_hwrite      ),
  .s3_req          (s3_req         ),
  .s4_haddr        (s4_haddr       ),
  .s4_hburst       (s4_hburst      ),
  .s4_hprot        (s4_hprot       ),
  .s4_hrdata       (s4_hrdata      ),
  .s4_hresp        (s4_hresp       ),
  .s4_hselx        (s4_hselx       ),
  .s4_hsize        (s4_hsize       ),
  .s4_htrans       (s4_htrans      ),
  .s4_hwdata       (s4_hwdata      ),
  .s4_hwrite       (s4_hwrite      ),
  .s4_req          (s4_req         ),
  .s5_haddr        (s5_haddr       ),
  .s5_hburst       (s5_hburst      ),
  .s5_hprot        (s5_hprot       ),
  .s5_hrdata       (s5_hrdata      ),
  .s5_hresp        (s5_hresp       ),
  .s5_hselx        (s5_hselx       ),
  .s5_hsize        (s5_hsize       ),
  .s5_htrans       (s5_htrans      ),
  .s5_hwdata       (s5_hwdata      ),
  .s5_hwrite       (s5_hwrite      ),
  .s5_req          (s5_req         ),
  .s6_haddr        (s6_haddr       ),
  .s6_hburst       (s6_hburst      ),
  .s6_hprot        (s6_hprot       ),
  .s6_hrdata       (s6_hrdata      ),
  .s6_hresp        (s6_hresp       ),
  .s6_hselx        (s6_hselx       ),
  .s6_hsize        (s6_hsize       ),
  .s6_htrans       (s6_htrans      ),
  .s6_hwdata       (s6_hwdata      ),
  .s6_hwrite       (s6_hwrite      ),
  .s6_req          (s6_req         ),
  .s7_haddr        (s7_haddr       ),
  .s7_hburst       (s7_hburst      ),
  .s7_hprot        (s7_hprot       ),
  .s7_hrdata       (s7_hrdata      ),
  .s7_hresp        (s7_hresp       ),
  .s7_hselx        (s7_hselx       ),
  .s7_hsize        (s7_hsize       ),
  .s7_htrans       (s7_htrans      ),
  .s7_hwdata       (s7_hwdata      ),
  .s7_hwrite       (s7_hwrite      ),
  .s7_req          (s7_req         ),
  .s8_haddr        (s8_haddr       ),
  .s8_hburst       (s8_hburst      ),
  .s8_hprot        (s8_hprot       ),
  .s8_hrdata       (s8_hrdata      ),
  .s8_hresp        (s8_hresp       ),
  .s8_hselx        (s8_hselx       ),
  .s8_hsize        (s8_hsize       ),
  .s8_htrans       (s8_htrans      ),
  .s8_hwdata       (s8_hwdata      ),
  .s8_hwrite       (s8_hwrite      ),
  .s8_req          (s8_req         ),
  .s9_haddr        (s9_haddr       ),
  .s9_hburst       (s9_hburst      ),
  .s9_hprot        (s9_hprot       ),
  .s9_hrdata       (s9_hrdata      ),
  .s9_hresp        (s9_hresp       ),
  .s9_hselx        (s9_hselx       ),
  .s9_hsize        (s9_hsize       ),
  .s9_htrans       (s9_htrans      ),
  .s9_hwdata       (s9_hwdata      ),
  .s9_hwrite       (s9_hwrite      ),
  .s9_req          (s9_req         )
);
ahb_matrix_7_12_arb  x_matrix_arb (
  .hclk            (hclk           ),
  .hresetn         (hresetn        ),
  .m0_latch_cmd    (m0_latch_cmd   ),
  .m0_nor_hready   (m0_nor_hready  ),
  .m0_s0_cmd_cur   (m0_s0_cmd_cur  ),
  .m0_s0_cmd_last  (m0_s0_cmd_last ),
  .m0_s0_data      (m0_s0_data     ),
  .m0_s0_req       (m0_s0_req      ),
  .m0_s10_cmd_cur  (m0_s10_cmd_cur ),
  .m0_s10_cmd_last (m0_s10_cmd_last),
  .m0_s10_data     (m0_s10_data    ),
  .m0_s10_req      (m0_s10_req     ),
  .m0_s11_cmd_cur  (m0_s11_cmd_cur ),
  .m0_s11_cmd_last (m0_s11_cmd_last),
  .m0_s11_data     (m0_s11_data    ),
  .m0_s11_req      (m0_s11_req     ),
  .m0_s1_cmd_cur   (m0_s1_cmd_cur  ),
  .m0_s1_cmd_last  (m0_s1_cmd_last ),
  .m0_s1_data      (m0_s1_data     ),
  .m0_s1_req       (m0_s1_req      ),
  .m0_s2_cmd_cur   (m0_s2_cmd_cur  ),
  .m0_s2_cmd_last  (m0_s2_cmd_last ),
  .m0_s2_data      (m0_s2_data     ),
  .m0_s2_req       (m0_s2_req      ),
  .m0_s3_cmd_cur   (m0_s3_cmd_cur  ),
  .m0_s3_cmd_last  (m0_s3_cmd_last ),
  .m0_s3_data      (m0_s3_data     ),
  .m0_s3_req       (m0_s3_req      ),
  .m0_s4_cmd_cur   (m0_s4_cmd_cur  ),
  .m0_s4_cmd_last  (m0_s4_cmd_last ),
  .m0_s4_data      (m0_s4_data     ),
  .m0_s4_req       (m0_s4_req      ),
  .m0_s5_cmd_cur   (m0_s5_cmd_cur  ),
  .m0_s5_cmd_last  (m0_s5_cmd_last ),
  .m0_s5_data      (m0_s5_data     ),
  .m0_s5_req       (m0_s5_req      ),
  .m0_s6_cmd_cur   (m0_s6_cmd_cur  ),
  .m0_s6_cmd_last  (m0_s6_cmd_last ),
  .m0_s6_data      (m0_s6_data     ),
  .m0_s6_req       (m0_s6_req      ),
  .m0_s7_cmd_cur   (m0_s7_cmd_cur  ),
  .m0_s7_cmd_last  (m0_s7_cmd_last ),
  .m0_s7_data      (m0_s7_data     ),
  .m0_s7_req       (m0_s7_req      ),
  .m0_s8_cmd_cur   (m0_s8_cmd_cur  ),
  .m0_s8_cmd_last  (m0_s8_cmd_last ),
  .m0_s8_data      (m0_s8_data     ),
  .m0_s8_req       (m0_s8_req      ),
  .m0_s9_cmd_cur   (m0_s9_cmd_cur  ),
  .m0_s9_cmd_last  (m0_s9_cmd_last ),
  .m0_s9_data      (m0_s9_data     ),
  .m0_s9_req       (m0_s9_req      ),
  .m1_latch_cmd    (m1_latch_cmd   ),
  .m1_nor_hready   (m1_nor_hready  ),
  .m1_s0_cmd_cur   (m1_s0_cmd_cur  ),
  .m1_s0_cmd_last  (m1_s0_cmd_last ),
  .m1_s0_data      (m1_s0_data     ),
  .m1_s0_req       (m1_s0_req      ),
  .m1_s10_cmd_cur  (m1_s10_cmd_cur ),
  .m1_s10_cmd_last (m1_s10_cmd_last),
  .m1_s10_data     (m1_s10_data    ),
  .m1_s10_req      (m1_s10_req     ),
  .m1_s11_cmd_cur  (m1_s11_cmd_cur ),
  .m1_s11_cmd_last (m1_s11_cmd_last),
  .m1_s11_data     (m1_s11_data    ),
  .m1_s11_req      (m1_s11_req     ),
  .m1_s1_cmd_cur   (m1_s1_cmd_cur  ),
  .m1_s1_cmd_last  (m1_s1_cmd_last ),
  .m1_s1_data      (m1_s1_data     ),
  .m1_s1_req       (m1_s1_req      ),
  .m1_s2_cmd_cur   (m1_s2_cmd_cur  ),
  .m1_s2_cmd_last  (m1_s2_cmd_last ),
  .m1_s2_data      (m1_s2_data     ),
  .m1_s2_req       (m1_s2_req      ),
  .m1_s3_cmd_cur   (m1_s3_cmd_cur  ),
  .m1_s3_cmd_last  (m1_s3_cmd_last ),
  .m1_s3_data      (m1_s3_data     ),
  .m1_s3_req       (m1_s3_req      ),
  .m1_s4_cmd_cur   (m1_s4_cmd_cur  ),
  .m1_s4_cmd_last  (m1_s4_cmd_last ),
  .m1_s4_data      (m1_s4_data     ),
  .m1_s4_req       (m1_s4_req      ),
  .m1_s5_cmd_cur   (m1_s5_cmd_cur  ),
  .m1_s5_cmd_last  (m1_s5_cmd_last ),
  .m1_s5_data      (m1_s5_data     ),
  .m1_s5_req       (m1_s5_req      ),
  .m1_s6_cmd_cur   (m1_s6_cmd_cur  ),
  .m1_s6_cmd_last  (m1_s6_cmd_last ),
  .m1_s6_data      (m1_s6_data     ),
  .m1_s6_req       (m1_s6_req      ),
  .m1_s7_cmd_cur   (m1_s7_cmd_cur  ),
  .m1_s7_cmd_last  (m1_s7_cmd_last ),
  .m1_s7_data      (m1_s7_data     ),
  .m1_s7_req       (m1_s7_req      ),
  .m1_s8_cmd_cur   (m1_s8_cmd_cur  ),
  .m1_s8_cmd_last  (m1_s8_cmd_last ),
  .m1_s8_data      (m1_s8_data     ),
  .m1_s8_req       (m1_s8_req      ),
  .m1_s9_cmd_cur   (m1_s9_cmd_cur  ),
  .m1_s9_cmd_last  (m1_s9_cmd_last ),
  .m1_s9_data      (m1_s9_data     ),
  .m1_s9_req       (m1_s9_req      ),
  .m2_latch_cmd    (m2_latch_cmd   ),
  .m2_nor_hready   (m2_nor_hready  ),
  .m2_s0_cmd_cur   (m2_s0_cmd_cur  ),
  .m2_s0_cmd_last  (m2_s0_cmd_last ),
  .m2_s0_data      (m2_s0_data     ),
  .m2_s0_req       (m2_s0_req      ),
  .m2_s10_cmd_cur  (m2_s10_cmd_cur ),
  .m2_s10_cmd_last (m2_s10_cmd_last),
  .m2_s10_data     (m2_s10_data    ),
  .m2_s10_req      (m2_s10_req     ),
  .m2_s11_cmd_cur  (m2_s11_cmd_cur ),
  .m2_s11_cmd_last (m2_s11_cmd_last),
  .m2_s11_data     (m2_s11_data    ),
  .m2_s11_req      (m2_s11_req     ),
  .m2_s1_cmd_cur   (m2_s1_cmd_cur  ),
  .m2_s1_cmd_last  (m2_s1_cmd_last ),
  .m2_s1_data      (m2_s1_data     ),
  .m2_s1_req       (m2_s1_req      ),
  .m2_s2_cmd_cur   (m2_s2_cmd_cur  ),
  .m2_s2_cmd_last  (m2_s2_cmd_last ),
  .m2_s2_data      (m2_s2_data     ),
  .m2_s2_req       (m2_s2_req      ),
  .m2_s3_cmd_cur   (m2_s3_cmd_cur  ),
  .m2_s3_cmd_last  (m2_s3_cmd_last ),
  .m2_s3_data      (m2_s3_data     ),
  .m2_s3_req       (m2_s3_req      ),
  .m2_s4_cmd_cur   (m2_s4_cmd_cur  ),
  .m2_s4_cmd_last  (m2_s4_cmd_last ),
  .m2_s4_data      (m2_s4_data     ),
  .m2_s4_req       (m2_s4_req      ),
  .m2_s5_cmd_cur   (m2_s5_cmd_cur  ),
  .m2_s5_cmd_last  (m2_s5_cmd_last ),
  .m2_s5_data      (m2_s5_data     ),
  .m2_s5_req       (m2_s5_req      ),
  .m2_s6_cmd_cur   (m2_s6_cmd_cur  ),
  .m2_s6_cmd_last  (m2_s6_cmd_last ),
  .m2_s6_data      (m2_s6_data     ),
  .m2_s6_req       (m2_s6_req      ),
  .m2_s7_cmd_cur   (m2_s7_cmd_cur  ),
  .m2_s7_cmd_last  (m2_s7_cmd_last ),
  .m2_s7_data      (m2_s7_data     ),
  .m2_s7_req       (m2_s7_req      ),
  .m2_s8_cmd_cur   (m2_s8_cmd_cur  ),
  .m2_s8_cmd_last  (m2_s8_cmd_last ),
  .m2_s8_data      (m2_s8_data     ),
  .m2_s8_req       (m2_s8_req      ),
  .m2_s9_cmd_cur   (m2_s9_cmd_cur  ),
  .m2_s9_cmd_last  (m2_s9_cmd_last ),
  .m2_s9_data      (m2_s9_data     ),
  .m2_s9_req       (m2_s9_req      ),
  .m3_latch_cmd    (m3_latch_cmd   ),
  .m3_nor_hready   (m3_nor_hready  ),
  .m3_s0_cmd_cur   (m3_s0_cmd_cur  ),
  .m3_s0_cmd_last  (m3_s0_cmd_last ),
  .m3_s0_data      (m3_s0_data     ),
  .m3_s0_req       (m3_s0_req      ),
  .m3_s10_cmd_cur  (m3_s10_cmd_cur ),
  .m3_s10_cmd_last (m3_s10_cmd_last),
  .m3_s10_data     (m3_s10_data    ),
  .m3_s10_req      (m3_s10_req     ),
  .m3_s11_cmd_cur  (m3_s11_cmd_cur ),
  .m3_s11_cmd_last (m3_s11_cmd_last),
  .m3_s11_data     (m3_s11_data    ),
  .m3_s11_req      (m3_s11_req     ),
  .m3_s1_cmd_cur   (m3_s1_cmd_cur  ),
  .m3_s1_cmd_last  (m3_s1_cmd_last ),
  .m3_s1_data      (m3_s1_data     ),
  .m3_s1_req       (m3_s1_req      ),
  .m3_s2_cmd_cur   (m3_s2_cmd_cur  ),
  .m3_s2_cmd_last  (m3_s2_cmd_last ),
  .m3_s2_data      (m3_s2_data     ),
  .m3_s2_req       (m3_s2_req      ),
  .m3_s3_cmd_cur   (m3_s3_cmd_cur  ),
  .m3_s3_cmd_last  (m3_s3_cmd_last ),
  .m3_s3_data      (m3_s3_data     ),
  .m3_s3_req       (m3_s3_req      ),
  .m3_s4_cmd_cur   (m3_s4_cmd_cur  ),
  .m3_s4_cmd_last  (m3_s4_cmd_last ),
  .m3_s4_data      (m3_s4_data     ),
  .m3_s4_req       (m3_s4_req      ),
  .m3_s5_cmd_cur   (m3_s5_cmd_cur  ),
  .m3_s5_cmd_last  (m3_s5_cmd_last ),
  .m3_s5_data      (m3_s5_data     ),
  .m3_s5_req       (m3_s5_req      ),
  .m3_s6_cmd_cur   (m3_s6_cmd_cur  ),
  .m3_s6_cmd_last  (m3_s6_cmd_last ),
  .m3_s6_data      (m3_s6_data     ),
  .m3_s6_req       (m3_s6_req      ),
  .m3_s7_cmd_cur   (m3_s7_cmd_cur  ),
  .m3_s7_cmd_last  (m3_s7_cmd_last ),
  .m3_s7_data      (m3_s7_data     ),
  .m3_s7_req       (m3_s7_req      ),
  .m3_s8_cmd_cur   (m3_s8_cmd_cur  ),
  .m3_s8_cmd_last  (m3_s8_cmd_last ),
  .m3_s8_data      (m3_s8_data     ),
  .m3_s8_req       (m3_s8_req      ),
  .m3_s9_cmd_cur   (m3_s9_cmd_cur  ),
  .m3_s9_cmd_last  (m3_s9_cmd_last ),
  .m3_s9_data      (m3_s9_data     ),
  .m3_s9_req       (m3_s9_req      ),
  .m4_latch_cmd    (m4_latch_cmd   ),
  .m4_nor_hready   (m4_nor_hready  ),
  .m4_s0_cmd_cur   (m4_s0_cmd_cur  ),
  .m4_s0_cmd_last  (m4_s0_cmd_last ),
  .m4_s0_data      (m4_s0_data     ),
  .m4_s0_req       (m4_s0_req      ),
  .m4_s10_cmd_cur  (m4_s10_cmd_cur ),
  .m4_s10_cmd_last (m4_s10_cmd_last),
  .m4_s10_data     (m4_s10_data    ),
  .m4_s10_req      (m4_s10_req     ),
  .m4_s11_cmd_cur  (m4_s11_cmd_cur ),
  .m4_s11_cmd_last (m4_s11_cmd_last),
  .m4_s11_data     (m4_s11_data    ),
  .m4_s11_req      (m4_s11_req     ),
  .m4_s1_cmd_cur   (m4_s1_cmd_cur  ),
  .m4_s1_cmd_last  (m4_s1_cmd_last ),
  .m4_s1_data      (m4_s1_data     ),
  .m4_s1_req       (m4_s1_req      ),
  .m4_s2_cmd_cur   (m4_s2_cmd_cur  ),
  .m4_s2_cmd_last  (m4_s2_cmd_last ),
  .m4_s2_data      (m4_s2_data     ),
  .m4_s2_req       (m4_s2_req      ),
  .m4_s3_cmd_cur   (m4_s3_cmd_cur  ),
  .m4_s3_cmd_last  (m4_s3_cmd_last ),
  .m4_s3_data      (m4_s3_data     ),
  .m4_s3_req       (m4_s3_req      ),
  .m4_s4_cmd_cur   (m4_s4_cmd_cur  ),
  .m4_s4_cmd_last  (m4_s4_cmd_last ),
  .m4_s4_data      (m4_s4_data     ),
  .m4_s4_req       (m4_s4_req      ),
  .m4_s5_cmd_cur   (m4_s5_cmd_cur  ),
  .m4_s5_cmd_last  (m4_s5_cmd_last ),
  .m4_s5_data      (m4_s5_data     ),
  .m4_s5_req       (m4_s5_req      ),
  .m4_s6_cmd_cur   (m4_s6_cmd_cur  ),
  .m4_s6_cmd_last  (m4_s6_cmd_last ),
  .m4_s6_data      (m4_s6_data     ),
  .m4_s6_req       (m4_s6_req      ),
  .m4_s7_cmd_cur   (m4_s7_cmd_cur  ),
  .m4_s7_cmd_last  (m4_s7_cmd_last ),
  .m4_s7_data      (m4_s7_data     ),
  .m4_s7_req       (m4_s7_req      ),
  .m4_s8_cmd_cur   (m4_s8_cmd_cur  ),
  .m4_s8_cmd_last  (m4_s8_cmd_last ),
  .m4_s8_data      (m4_s8_data     ),
  .m4_s8_req       (m4_s8_req      ),
  .m4_s9_cmd_cur   (m4_s9_cmd_cur  ),
  .m4_s9_cmd_last  (m4_s9_cmd_last ),
  .m4_s9_data      (m4_s9_data     ),
  .m4_s9_req       (m4_s9_req      ),
  .m5_latch_cmd    (m5_latch_cmd   ),
  .m5_nor_hready   (m5_nor_hready  ),
  .m5_s0_cmd_cur   (m5_s0_cmd_cur  ),
  .m5_s0_cmd_last  (m5_s0_cmd_last ),
  .m5_s0_data      (m5_s0_data     ),
  .m5_s0_req       (m5_s0_req      ),
  .m5_s10_cmd_cur  (m5_s10_cmd_cur ),
  .m5_s10_cmd_last (m5_s10_cmd_last),
  .m5_s10_data     (m5_s10_data    ),
  .m5_s10_req      (m5_s10_req     ),
  .m5_s11_cmd_cur  (m5_s11_cmd_cur ),
  .m5_s11_cmd_last (m5_s11_cmd_last),
  .m5_s11_data     (m5_s11_data    ),
  .m5_s11_req      (m5_s11_req     ),
  .m5_s1_cmd_cur   (m5_s1_cmd_cur  ),
  .m5_s1_cmd_last  (m5_s1_cmd_last ),
  .m5_s1_data      (m5_s1_data     ),
  .m5_s1_req       (m5_s1_req      ),
  .m5_s2_cmd_cur   (m5_s2_cmd_cur  ),
  .m5_s2_cmd_last  (m5_s2_cmd_last ),
  .m5_s2_data      (m5_s2_data     ),
  .m5_s2_req       (m5_s2_req      ),
  .m5_s3_cmd_cur   (m5_s3_cmd_cur  ),
  .m5_s3_cmd_last  (m5_s3_cmd_last ),
  .m5_s3_data      (m5_s3_data     ),
  .m5_s3_req       (m5_s3_req      ),
  .m5_s4_cmd_cur   (m5_s4_cmd_cur  ),
  .m5_s4_cmd_last  (m5_s4_cmd_last ),
  .m5_s4_data      (m5_s4_data     ),
  .m5_s4_req       (m5_s4_req      ),
  .m5_s5_cmd_cur   (m5_s5_cmd_cur  ),
  .m5_s5_cmd_last  (m5_s5_cmd_last ),
  .m5_s5_data      (m5_s5_data     ),
  .m5_s5_req       (m5_s5_req      ),
  .m5_s6_cmd_cur   (m5_s6_cmd_cur  ),
  .m5_s6_cmd_last  (m5_s6_cmd_last ),
  .m5_s6_data      (m5_s6_data     ),
  .m5_s6_req       (m5_s6_req      ),
  .m5_s7_cmd_cur   (m5_s7_cmd_cur  ),
  .m5_s7_cmd_last  (m5_s7_cmd_last ),
  .m5_s7_data      (m5_s7_data     ),
  .m5_s7_req       (m5_s7_req      ),
  .m5_s8_cmd_cur   (m5_s8_cmd_cur  ),
  .m5_s8_cmd_last  (m5_s8_cmd_last ),
  .m5_s8_data      (m5_s8_data     ),
  .m5_s8_req       (m5_s8_req      ),
  .m5_s9_cmd_cur   (m5_s9_cmd_cur  ),
  .m5_s9_cmd_last  (m5_s9_cmd_last ),
  .m5_s9_data      (m5_s9_data     ),
  .m5_s9_req       (m5_s9_req      ),
  .m6_latch_cmd    (m6_latch_cmd   ),
  .m6_nor_hready   (m6_nor_hready  ),
  .m6_s0_cmd_cur   (m6_s0_cmd_cur  ),
  .m6_s0_cmd_last  (m6_s0_cmd_last ),
  .m6_s0_data      (m6_s0_data     ),
  .m6_s0_req       (m6_s0_req      ),
  .m6_s10_cmd_cur  (m6_s10_cmd_cur ),
  .m6_s10_cmd_last (m6_s10_cmd_last),
  .m6_s10_data     (m6_s10_data    ),
  .m6_s10_req      (m6_s10_req     ),
  .m6_s11_cmd_cur  (m6_s11_cmd_cur ),
  .m6_s11_cmd_last (m6_s11_cmd_last),
  .m6_s11_data     (m6_s11_data    ),
  .m6_s11_req      (m6_s11_req     ),
  .m6_s1_cmd_cur   (m6_s1_cmd_cur  ),
  .m6_s1_cmd_last  (m6_s1_cmd_last ),
  .m6_s1_data      (m6_s1_data     ),
  .m6_s1_req       (m6_s1_req      ),
  .m6_s2_cmd_cur   (m6_s2_cmd_cur  ),
  .m6_s2_cmd_last  (m6_s2_cmd_last ),
  .m6_s2_data      (m6_s2_data     ),
  .m6_s2_req       (m6_s2_req      ),
  .m6_s3_cmd_cur   (m6_s3_cmd_cur  ),
  .m6_s3_cmd_last  (m6_s3_cmd_last ),
  .m6_s3_data      (m6_s3_data     ),
  .m6_s3_req       (m6_s3_req      ),
  .m6_s4_cmd_cur   (m6_s4_cmd_cur  ),
  .m6_s4_cmd_last  (m6_s4_cmd_last ),
  .m6_s4_data      (m6_s4_data     ),
  .m6_s4_req       (m6_s4_req      ),
  .m6_s5_cmd_cur   (m6_s5_cmd_cur  ),
  .m6_s5_cmd_last  (m6_s5_cmd_last ),
  .m6_s5_data      (m6_s5_data     ),
  .m6_s5_req       (m6_s5_req      ),
  .m6_s6_cmd_cur   (m6_s6_cmd_cur  ),
  .m6_s6_cmd_last  (m6_s6_cmd_last ),
  .m6_s6_data      (m6_s6_data     ),
  .m6_s6_req       (m6_s6_req      ),
  .m6_s7_cmd_cur   (m6_s7_cmd_cur  ),
  .m6_s7_cmd_last  (m6_s7_cmd_last ),
  .m6_s7_data      (m6_s7_data     ),
  .m6_s7_req       (m6_s7_req      ),
  .m6_s8_cmd_cur   (m6_s8_cmd_cur  ),
  .m6_s8_cmd_last  (m6_s8_cmd_last ),
  .m6_s8_data      (m6_s8_data     ),
  .m6_s8_req       (m6_s8_req      ),
  .m6_s9_cmd_cur   (m6_s9_cmd_cur  ),
  .m6_s9_cmd_last  (m6_s9_cmd_last ),
  .m6_s9_data      (m6_s9_data     ),
  .m6_s9_req       (m6_s9_req      ),
  .s0_hready       (s0_hready      ),
  .s0_req          (s0_req         ),
  .s10_hready      (s10_hready     ),
  .s10_req         (s10_req        ),
  .s11_hready      (s11_hready     ),
  .s11_req         (s11_req        ),
  .s1_hready       (s1_hready      ),
  .s1_req          (s1_req         ),
  .s2_hready       (s2_hready      ),
  .s2_req          (s2_req         ),
  .s3_hready       (s3_hready      ),
  .s3_req          (s3_req         ),
  .s4_hready       (s4_hready      ),
  .s4_req          (s4_req         ),
  .s5_hready       (s5_hready      ),
  .s5_req          (s5_req         ),
  .s6_hready       (s6_hready      ),
  .s6_req          (s6_req         ),
  .s7_hready       (s7_hready      ),
  .s7_req          (s7_req         ),
  .s8_hready       (s8_hready      ),
  .s8_req          (s8_req         ),
  .s9_hready       (s9_hready      ),
  .s9_req          (s9_req         )
);
endmodule
